VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu8bit
  CLASS BLOCK ;
  FOREIGN alu8bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.445 BY 91.165 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 79.120 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 79.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 74.760 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.730 74.760 78.330 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 76.445 54.440 80.445 55.040 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 76.445 30.640 80.445 31.240 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 87.165 22.910 91.165 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 87.165 67.990 91.165 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 87.165 77.650 91.165 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 87.165 58.330 91.165 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 76.445 6.840 80.445 7.440 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 87.165 0.370 91.165 ;
    END
  END b[7]
  PIN carry
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END carry
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 87.165 45.450 91.165 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END opcode[1]
  PIN opcode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 87.165 13.250 91.165 ;
    END
  END opcode[2]
  PIN opcode[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 76.445 20.440 80.445 21.040 ;
    END
  END opcode[3]
  PIN result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END result[0]
  PIN result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 76.445 68.040 80.445 68.640 ;
    END
  END result[1]
  PIN result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 76.445 78.240 80.445 78.840 ;
    END
  END result[2]
  PIN result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 87.165 35.790 91.165 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END result[7]
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 76.445 44.240 80.445 44.840 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.520 78.965 ;
      LAYER met1 ;
        RECT 0.070 10.640 77.670 79.120 ;
      LAYER met2 ;
        RECT 0.650 86.885 12.690 87.165 ;
        RECT 13.530 86.885 22.350 87.165 ;
        RECT 23.190 86.885 35.230 87.165 ;
        RECT 36.070 86.885 44.890 87.165 ;
        RECT 45.730 86.885 57.770 87.165 ;
        RECT 58.610 86.885 67.430 87.165 ;
        RECT 68.270 86.885 77.090 87.165 ;
        RECT 0.100 4.280 77.640 86.885 ;
        RECT 0.650 4.000 9.470 4.280 ;
        RECT 10.310 4.000 19.130 4.280 ;
        RECT 19.970 4.000 32.010 4.280 ;
        RECT 32.850 4.000 41.670 4.280 ;
        RECT 42.510 4.000 54.550 4.280 ;
        RECT 55.390 4.000 64.210 4.280 ;
        RECT 65.050 4.000 77.090 4.280 ;
      LAYER met3 ;
        RECT 4.400 81.240 76.445 82.105 ;
        RECT 4.000 79.240 76.445 81.240 ;
        RECT 4.000 77.840 76.045 79.240 ;
        RECT 4.000 69.040 76.445 77.840 ;
        RECT 4.400 67.640 76.045 69.040 ;
        RECT 4.000 58.840 76.445 67.640 ;
        RECT 4.400 57.440 76.445 58.840 ;
        RECT 4.000 55.440 76.445 57.440 ;
        RECT 4.000 54.040 76.045 55.440 ;
        RECT 4.000 45.240 76.445 54.040 ;
        RECT 4.400 43.840 76.045 45.240 ;
        RECT 4.000 35.040 76.445 43.840 ;
        RECT 4.400 33.640 76.445 35.040 ;
        RECT 4.000 31.640 76.445 33.640 ;
        RECT 4.000 30.240 76.045 31.640 ;
        RECT 4.000 21.440 76.445 30.240 ;
        RECT 4.400 20.040 76.045 21.440 ;
        RECT 4.000 11.240 76.445 20.040 ;
        RECT 4.400 9.840 76.445 11.240 ;
        RECT 4.000 7.840 76.445 9.840 ;
        RECT 4.000 6.975 76.045 7.840 ;
      LAYER met4 ;
        RECT 34.335 19.895 34.665 41.985 ;
  END
END alu8bit
END LIBRARY

