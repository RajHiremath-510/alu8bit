magic
tech sky130A
magscale 1 2
timestamp 1755626710
<< checkpaint >>
rect -3932 -3932 20021 22165
<< viali >>
rect 1501 15657 1535 15691
rect 7297 15657 7331 15691
rect 14289 15657 14323 15691
rect 1961 15453 1995 15487
rect 2697 15453 2731 15487
rect 4629 15453 4663 15487
rect 9321 15453 9355 15487
rect 11805 15453 11839 15487
rect 13921 15453 13955 15487
rect 1777 15385 1811 15419
rect 7573 15385 7607 15419
rect 14197 15385 14231 15419
rect 2145 15317 2179 15351
rect 2881 15317 2915 15351
rect 4813 15317 4847 15351
rect 9137 15317 9171 15351
rect 11897 15317 11931 15351
rect 13737 15317 13771 15351
rect 14473 15113 14507 15147
rect 14197 14977 14231 15011
rect 1409 13889 1443 13923
rect 7297 13889 7331 13923
rect 14197 13889 14231 13923
rect 1685 13821 1719 13855
rect 7389 13821 7423 13855
rect 14473 13821 14507 13855
rect 7665 13753 7699 13787
rect 4537 13481 4571 13515
rect 5089 13481 5123 13515
rect 9689 13413 9723 13447
rect 5273 13345 5307 13379
rect 5457 13345 5491 13379
rect 5917 13345 5951 13379
rect 8585 13345 8619 13379
rect 9137 13345 9171 13379
rect 9965 13345 9999 13379
rect 10057 13345 10091 13379
rect 4261 13277 4295 13311
rect 4813 13277 4847 13311
rect 5549 13277 5583 13311
rect 6561 13277 6595 13311
rect 7481 13277 7515 13311
rect 8309 13277 8343 13311
rect 8401 13277 8435 13311
rect 8493 13277 8527 13311
rect 9229 13277 9263 13311
rect 9873 13277 9907 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 10517 13277 10551 13311
rect 10701 13277 10735 13311
rect 10793 13277 10827 13311
rect 8033 13209 8067 13243
rect 4721 13141 4755 13175
rect 8125 13141 8159 13175
rect 9597 13141 9631 13175
rect 10425 13141 10459 13175
rect 5181 12937 5215 12971
rect 7389 12937 7423 12971
rect 8854 12937 8888 12971
rect 10425 12937 10459 12971
rect 5089 12869 5123 12903
rect 5273 12869 5307 12903
rect 8953 12869 8987 12903
rect 11529 12869 11563 12903
rect 4353 12801 4387 12835
rect 4445 12801 4479 12835
rect 4629 12801 4663 12835
rect 4997 12801 5031 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7665 12801 7699 12835
rect 7757 12801 7791 12835
rect 7941 12801 7975 12835
rect 8677 12801 8711 12835
rect 8769 12801 8803 12835
rect 10885 12801 10919 12835
rect 12449 12801 12483 12835
rect 13369 12801 13403 12835
rect 8309 12665 8343 12699
rect 10609 12665 10643 12699
rect 4813 12597 4847 12631
rect 6101 12189 6135 12223
rect 6285 12189 6319 12223
rect 6285 12053 6319 12087
rect 4721 11849 4755 11883
rect 5549 11849 5583 11883
rect 9505 11849 9539 11883
rect 10241 11849 10275 11883
rect 11069 11849 11103 11883
rect 1777 11781 1811 11815
rect 5181 11781 5215 11815
rect 7757 11781 7791 11815
rect 9873 11781 9907 11815
rect 9965 11781 9999 11815
rect 10609 11781 10643 11815
rect 1409 11713 1443 11747
rect 3893 11713 3927 11747
rect 4629 11713 4663 11747
rect 5365 11713 5399 11747
rect 5549 11713 5583 11747
rect 5641 11713 5675 11747
rect 5733 11713 5767 11747
rect 5917 11713 5951 11747
rect 6009 11713 6043 11747
rect 6653 11713 6687 11747
rect 6745 11713 6779 11747
rect 7941 11713 7975 11747
rect 8217 11713 8251 11747
rect 8309 11713 8343 11747
rect 9137 11713 9171 11747
rect 9597 11713 9631 11747
rect 9745 11713 9779 11747
rect 10062 11713 10096 11747
rect 10793 11713 10827 11747
rect 10977 11713 11011 11747
rect 11253 11713 11287 11747
rect 3985 11645 4019 11679
rect 6377 11645 6411 11679
rect 6561 11645 6595 11679
rect 6837 11645 6871 11679
rect 8033 11645 8067 11679
rect 9229 11645 9263 11679
rect 4813 11577 4847 11611
rect 6193 11577 6227 11611
rect 7573 11509 7607 11543
rect 8125 11509 8159 11543
rect 5089 11305 5123 11339
rect 6469 11305 6503 11339
rect 9781 11305 9815 11339
rect 10885 11305 10919 11339
rect 11345 11305 11379 11339
rect 8401 11237 8435 11271
rect 4629 11169 4663 11203
rect 14289 11169 14323 11203
rect 4537 11101 4571 11135
rect 4813 11101 4847 11135
rect 4905 11101 4939 11135
rect 5181 11101 5215 11135
rect 5365 11101 5399 11135
rect 6101 11101 6135 11135
rect 7297 11101 7331 11135
rect 7573 11101 7607 11135
rect 7849 11101 7883 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 8217 11101 8251 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 11069 11101 11103 11135
rect 11161 11101 11195 11135
rect 11437 11101 11471 11135
rect 14565 11101 14599 11135
rect 5273 11033 5307 11067
rect 6285 11033 6319 11067
rect 7389 11033 7423 11067
rect 7757 11033 7791 11067
rect 9137 11033 9171 11067
rect 4629 10761 4663 10795
rect 8059 10761 8093 10795
rect 11161 10761 11195 10795
rect 7849 10693 7883 10727
rect 4169 10625 4203 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 4721 10625 4755 10659
rect 11069 10625 11103 10659
rect 11253 10625 11287 10659
rect 3985 10557 4019 10591
rect 8033 10421 8067 10455
rect 8217 10421 8251 10455
rect 8493 10217 8527 10251
rect 9873 10217 9907 10251
rect 10149 10217 10183 10251
rect 11069 10217 11103 10251
rect 6285 10149 6319 10183
rect 6377 10081 6411 10115
rect 6745 10081 6779 10115
rect 6837 10081 6871 10115
rect 8309 10081 8343 10115
rect 4077 10013 4111 10047
rect 4225 10013 4259 10047
rect 4445 10013 4479 10047
rect 4583 10013 4617 10047
rect 5641 10013 5675 10047
rect 5734 10013 5768 10047
rect 6147 10013 6181 10047
rect 6561 10013 6595 10047
rect 7021 10013 7055 10047
rect 7193 10013 7227 10047
rect 7300 10013 7334 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 8585 10013 8619 10047
rect 9229 10013 9263 10047
rect 9377 10013 9411 10047
rect 9735 10013 9769 10047
rect 10425 10013 10459 10047
rect 10517 10013 10551 10047
rect 10609 10013 10643 10047
rect 10793 10013 10827 10047
rect 11253 10013 11287 10047
rect 11437 10013 11471 10047
rect 4353 9945 4387 9979
rect 5917 9945 5951 9979
rect 6009 9945 6043 9979
rect 9505 9945 9539 9979
rect 9597 9945 9631 9979
rect 4721 9877 4755 9911
rect 7757 9877 7791 9911
rect 8033 9877 8067 9911
rect 3709 9673 3743 9707
rect 7849 9673 7883 9707
rect 9229 9673 9263 9707
rect 10149 9673 10183 9707
rect 4261 9605 4295 9639
rect 6653 9605 6687 9639
rect 9965 9605 9999 9639
rect 3985 9537 4019 9571
rect 4353 9537 4387 9571
rect 6469 9537 6503 9571
rect 6745 9537 6779 9571
rect 7481 9537 7515 9571
rect 9505 9537 9539 9571
rect 10149 9537 10183 9571
rect 10241 9537 10275 9571
rect 10333 9537 10367 9571
rect 10517 9537 10551 9571
rect 11713 9537 11747 9571
rect 11897 9537 11931 9571
rect 3893 9469 3927 9503
rect 9413 9469 9447 9503
rect 9781 9469 9815 9503
rect 9873 9469 9907 9503
rect 11989 9469 12023 9503
rect 6745 9401 6779 9435
rect 8033 9401 8067 9435
rect 7849 9333 7883 9367
rect 10333 9333 10367 9367
rect 11529 9333 11563 9367
rect 7711 9129 7745 9163
rect 10885 9129 10919 9163
rect 11529 9129 11563 9163
rect 7849 9061 7883 9095
rect 11069 9061 11103 9095
rect 3985 8993 4019 9027
rect 5365 8993 5399 9027
rect 7941 8993 7975 9027
rect 1777 8925 1811 8959
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 4593 8925 4627 8959
rect 4721 8925 4755 8959
rect 4951 8925 4985 8959
rect 5273 8925 5307 8959
rect 5549 8925 5583 8959
rect 5641 8925 5675 8959
rect 6653 8925 6687 8959
rect 7573 8925 7607 8959
rect 8309 8925 8343 8959
rect 9045 8925 9079 8959
rect 9413 8925 9447 8959
rect 9689 8925 9723 8959
rect 10149 8925 10183 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 12817 8925 12851 8959
rect 13185 8925 13219 8959
rect 10931 8891 10965 8925
rect 1409 8857 1443 8891
rect 4813 8857 4847 8891
rect 10701 8857 10735 8891
rect 11805 8857 11839 8891
rect 4353 8789 4387 8823
rect 5089 8789 5123 8823
rect 5825 8789 5859 8823
rect 6745 8789 6779 8823
rect 10333 8789 10367 8823
rect 11161 8789 11195 8823
rect 12173 8789 12207 8823
rect 4169 8585 4203 8619
rect 4905 8585 4939 8619
rect 5273 8585 5307 8619
rect 6653 8585 6687 8619
rect 7481 8585 7515 8619
rect 8953 8585 8987 8619
rect 11529 8585 11563 8619
rect 3525 8517 3559 8551
rect 9229 8517 9263 8551
rect 14473 8517 14507 8551
rect 4077 8449 4111 8483
rect 4261 8449 4295 8483
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 6837 8449 6871 8483
rect 7113 8449 7147 8483
rect 7573 8449 7607 8483
rect 7665 8449 7699 8483
rect 9137 8449 9171 8483
rect 9321 8449 9355 8483
rect 9505 8449 9539 8483
rect 9597 8449 9631 8483
rect 10149 8449 10183 8483
rect 10241 8449 10275 8483
rect 10425 8449 10459 8483
rect 10527 8455 10561 8489
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 12081 8449 12115 8483
rect 13921 8449 13955 8483
rect 7021 8381 7055 8415
rect 7205 8381 7239 8415
rect 7389 8381 7423 8415
rect 7297 8313 7331 8347
rect 7849 8313 7883 8347
rect 9965 8313 9999 8347
rect 11989 8313 12023 8347
rect 3433 8245 3467 8279
rect 5089 8245 5123 8279
rect 5273 8245 5307 8279
rect 6561 8041 6595 8075
rect 9413 8041 9447 8075
rect 4353 7973 4387 8007
rect 4445 7905 4479 7939
rect 8125 7905 8159 7939
rect 8217 7905 8251 7939
rect 8309 7905 8343 7939
rect 13093 7905 13127 7939
rect 2973 7837 3007 7871
rect 3893 7837 3927 7871
rect 3985 7837 4019 7871
rect 6469 7837 6503 7871
rect 6653 7837 6687 7871
rect 7021 7837 7055 7871
rect 8401 7837 8435 7871
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 9873 7837 9907 7871
rect 2789 7769 2823 7803
rect 12265 7769 12299 7803
rect 4721 7701 4755 7735
rect 6837 7701 6871 7735
rect 7941 7701 7975 7735
rect 8585 7497 8619 7531
rect 8769 7497 8803 7531
rect 9505 7497 9539 7531
rect 2053 7429 2087 7463
rect 3525 7429 3559 7463
rect 4077 7429 4111 7463
rect 6469 7429 6503 7463
rect 8125 7429 8159 7463
rect 11805 7429 11839 7463
rect 11897 7429 11931 7463
rect 1501 7361 1535 7395
rect 3065 7361 3099 7395
rect 3617 7361 3651 7395
rect 4261 7361 4295 7395
rect 6745 7361 6779 7395
rect 8677 7361 8711 7395
rect 8953 7361 8987 7395
rect 9873 7361 9907 7395
rect 11713 7361 11747 7395
rect 12081 7361 12115 7395
rect 3985 7293 4019 7327
rect 6653 7293 6687 7327
rect 9965 7293 9999 7327
rect 8493 7225 8527 7259
rect 9137 7225 9171 7259
rect 4445 7157 4479 7191
rect 6745 7157 6779 7191
rect 6929 7157 6963 7191
rect 10149 7157 10183 7191
rect 11529 7157 11563 7191
rect 4169 6953 4203 6987
rect 4353 6953 4387 6987
rect 4997 6953 5031 6987
rect 5181 6953 5215 6987
rect 5825 6953 5859 6987
rect 3525 6885 3559 6919
rect 6193 6885 6227 6919
rect 10609 6885 10643 6919
rect 3801 6817 3835 6851
rect 4629 6817 4663 6851
rect 8953 6817 8987 6851
rect 9597 6817 9631 6851
rect 9781 6817 9815 6851
rect 12725 6817 12759 6851
rect 12909 6817 12943 6851
rect 2973 6749 3007 6783
rect 3157 6749 3191 6783
rect 3341 6749 3375 6783
rect 5733 6749 5767 6783
rect 5825 6749 5859 6783
rect 6745 6749 6779 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 9505 6749 9539 6783
rect 9873 6749 9907 6783
rect 10057 6749 10091 6783
rect 10333 6749 10367 6783
rect 10425 6749 10459 6783
rect 10701 6749 10735 6783
rect 10885 6749 10919 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 11713 6749 11747 6783
rect 11805 6749 11839 6783
rect 11897 6749 11931 6783
rect 12633 6749 12667 6783
rect 13093 6749 13127 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 3065 6681 3099 6715
rect 4169 6681 4203 6715
rect 4997 6681 5031 6715
rect 5365 6681 5399 6715
rect 6193 6681 6227 6715
rect 9965 6681 9999 6715
rect 10609 6681 10643 6715
rect 6009 6613 6043 6647
rect 6653 6613 6687 6647
rect 6929 6613 6963 6647
rect 9321 6613 9355 6647
rect 9781 6613 9815 6647
rect 12173 6613 12207 6647
rect 12265 6613 12299 6647
rect 3801 6409 3835 6443
rect 4813 6409 4847 6443
rect 4997 6409 5031 6443
rect 7573 6409 7607 6443
rect 10609 6409 10643 6443
rect 12909 6409 12943 6443
rect 2789 6341 2823 6375
rect 4629 6341 4663 6375
rect 3249 6273 3283 6307
rect 3525 6273 3559 6307
rect 4261 6273 4295 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 7021 6273 7055 6307
rect 7113 6273 7147 6307
rect 8125 6273 8159 6307
rect 8585 6273 8619 6307
rect 8861 6273 8895 6307
rect 8953 6273 8987 6307
rect 9137 6273 9171 6307
rect 9229 6273 9263 6307
rect 9321 6273 9355 6307
rect 10425 6273 10459 6307
rect 10609 6273 10643 6307
rect 12817 6273 12851 6307
rect 14473 6273 14507 6307
rect 3157 6205 3191 6239
rect 3893 6205 3927 6239
rect 3985 6205 4019 6239
rect 7849 6205 7883 6239
rect 9781 6137 9815 6171
rect 2881 6069 2915 6103
rect 3433 6069 3467 6103
rect 4813 6069 4847 6103
rect 8677 6069 8711 6103
rect 9413 6069 9447 6103
rect 14381 6069 14415 6103
rect 3433 5865 3467 5899
rect 5365 5865 5399 5899
rect 7021 5865 7055 5899
rect 7941 5865 7975 5899
rect 8125 5865 8159 5899
rect 11161 5865 11195 5899
rect 12449 5865 12483 5899
rect 5549 5729 5583 5763
rect 6837 5729 6871 5763
rect 8033 5729 8067 5763
rect 3801 5661 3835 5695
rect 5089 5661 5123 5695
rect 6561 5661 6595 5695
rect 6653 5661 6687 5695
rect 6745 5661 6779 5695
rect 8254 5661 8288 5695
rect 11321 5661 11355 5695
rect 11713 5661 11747 5695
rect 12541 5661 12575 5695
rect 3525 5593 3559 5627
rect 8401 5593 8435 5627
rect 11437 5593 11471 5627
rect 11529 5593 11563 5627
rect 12725 5593 12759 5627
rect 3985 5525 4019 5559
rect 5549 5321 5583 5355
rect 8125 5321 8159 5355
rect 12357 5321 12391 5355
rect 13369 5321 13403 5355
rect 5365 5253 5399 5287
rect 6469 5253 6503 5287
rect 11253 5253 11287 5287
rect 4721 5185 4755 5219
rect 4813 5185 4847 5219
rect 5181 5185 5215 5219
rect 5641 5185 5675 5219
rect 5825 5185 5859 5219
rect 6745 5185 6779 5219
rect 6837 5185 6871 5219
rect 7941 5185 7975 5219
rect 8033 5185 8067 5219
rect 9597 5185 9631 5219
rect 10149 5185 10183 5219
rect 10425 5185 10459 5219
rect 10517 5185 10551 5219
rect 10885 5185 10919 5219
rect 12265 5185 12299 5219
rect 12449 5185 12483 5219
rect 13001 5185 13035 5219
rect 13093 5185 13127 5219
rect 13185 5185 13219 5219
rect 13461 5185 13495 5219
rect 4905 5117 4939 5151
rect 4997 5117 5031 5151
rect 6377 5117 6411 5151
rect 8309 5117 8343 5151
rect 9689 5117 9723 5151
rect 10057 5117 10091 5151
rect 10333 5117 10367 5151
rect 10793 5117 10827 5151
rect 11161 5117 11195 5151
rect 10149 5049 10183 5083
rect 4537 4981 4571 5015
rect 5641 4981 5675 5015
rect 7021 4981 7055 5015
rect 8033 4981 8067 5015
rect 9413 4981 9447 5015
rect 10609 4981 10643 5015
rect 12725 4981 12759 5015
rect 13093 4981 13127 5015
rect 13185 4981 13219 5015
rect 6653 4777 6687 4811
rect 7113 4777 7147 4811
rect 11253 4777 11287 4811
rect 12265 4777 12299 4811
rect 14381 4777 14415 4811
rect 7849 4709 7883 4743
rect 12357 4709 12391 4743
rect 6469 4641 6503 4675
rect 8125 4641 8159 4675
rect 8217 4641 8251 4675
rect 1409 4573 1443 4607
rect 4997 4573 5031 4607
rect 5181 4573 5215 4607
rect 6285 4573 6319 4607
rect 6653 4573 6687 4607
rect 6745 4573 6779 4607
rect 6929 4573 6963 4607
rect 8033 4573 8067 4607
rect 8309 4573 8343 4607
rect 9597 4573 9631 4607
rect 9689 4573 9723 4607
rect 9858 4573 9892 4607
rect 9965 4573 9999 4607
rect 11437 4573 11471 4607
rect 11529 4573 11563 4607
rect 12081 4573 12115 4607
rect 12725 4573 12759 4607
rect 14565 4573 14599 4607
rect 11897 4505 11931 4539
rect 1593 4437 1627 4471
rect 5181 4437 5215 4471
rect 6377 4437 6411 4471
rect 9413 4437 9447 4471
rect 11713 4437 11747 4471
rect 8953 4233 8987 4267
rect 5089 4165 5123 4199
rect 4721 4097 4755 4131
rect 4814 4097 4848 4131
rect 4997 4097 5031 4131
rect 5227 4097 5261 4131
rect 5457 4097 5491 4131
rect 5641 4097 5675 4131
rect 8125 4097 8159 4131
rect 9137 4097 9171 4131
rect 9321 4097 9355 4131
rect 9873 4097 9907 4131
rect 9965 4097 9999 4131
rect 10149 4097 10183 4131
rect 10241 4097 10275 4131
rect 11989 4097 12023 4131
rect 8217 4029 8251 4063
rect 8309 4029 8343 4063
rect 8401 4029 8435 4063
rect 9229 4029 9263 4063
rect 9413 4029 9447 4063
rect 9689 4029 9723 4063
rect 11529 3961 11563 3995
rect 5365 3893 5399 3927
rect 5549 3893 5583 3927
rect 7941 3893 7975 3927
rect 11713 3893 11747 3927
rect 7849 3689 7883 3723
rect 8217 3689 8251 3723
rect 9965 3689 9999 3723
rect 10241 3689 10275 3723
rect 6193 3621 6227 3655
rect 12081 3621 12115 3655
rect 5917 3553 5951 3587
rect 8125 3553 8159 3587
rect 10885 3553 10919 3587
rect 6101 3485 6135 3519
rect 6377 3485 6411 3519
rect 6469 3485 6503 3519
rect 8217 3485 8251 3519
rect 9781 3485 9815 3519
rect 10425 3485 10459 3519
rect 10609 3485 10643 3519
rect 6193 3417 6227 3451
rect 9597 3417 9631 3451
rect 10517 3417 10551 3451
rect 10727 3417 10761 3451
rect 11713 3417 11747 3451
rect 12173 3349 12207 3383
rect 6009 3145 6043 3179
rect 6469 3145 6503 3179
rect 9413 3145 9447 3179
rect 10149 3145 10183 3179
rect 12081 3145 12115 3179
rect 8953 3077 8987 3111
rect 10057 3077 10091 3111
rect 4997 3009 5031 3043
rect 5181 3009 5215 3043
rect 5273 3009 5307 3043
rect 5457 3009 5491 3043
rect 5549 3009 5583 3043
rect 5733 3009 5767 3043
rect 5825 3009 5859 3043
rect 6653 3009 6687 3043
rect 6929 3009 6963 3043
rect 7757 3009 7791 3043
rect 7849 3009 7883 3043
rect 7941 3009 7975 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 8769 3009 8803 3043
rect 9873 3009 9907 3043
rect 10333 3009 10367 3043
rect 10517 3009 10551 3043
rect 10617 3009 10651 3043
rect 10793 3009 10827 3043
rect 11069 3009 11103 3043
rect 11529 3009 11563 3043
rect 11805 3009 11839 3043
rect 11897 3009 11931 3043
rect 6745 2941 6779 2975
rect 6837 2941 6871 2975
rect 9689 2941 9723 2975
rect 4997 2873 5031 2907
rect 7481 2873 7515 2907
rect 8217 2873 8251 2907
rect 9229 2873 9263 2907
rect 10701 2873 10735 2907
rect 5457 2805 5491 2839
rect 5825 2805 5859 2839
rect 8677 2805 8711 2839
rect 10977 2805 11011 2839
rect 11621 2805 11655 2839
rect 2145 2601 2179 2635
rect 2513 2601 2547 2635
rect 4169 2601 4203 2635
rect 7665 2601 7699 2635
rect 11069 2601 11103 2635
rect 1777 2533 1811 2567
rect 7757 2533 7791 2567
rect 8125 2465 8159 2499
rect 8953 2465 8987 2499
rect 13277 2465 13311 2499
rect 2329 2397 2363 2431
rect 3985 2397 4019 2431
rect 6745 2397 6779 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 11253 2397 11287 2431
rect 12817 2397 12851 2431
rect 13093 2397 13127 2431
rect 13829 2397 13863 2431
rect 14197 2397 14231 2431
rect 1501 2329 1535 2363
rect 2053 2329 2087 2363
rect 8677 2329 8711 2363
rect 14565 2329 14599 2363
rect 6469 2261 6503 2295
rect 8401 2261 8435 2295
<< metal1 >>
rect 1104 15802 14904 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 14214 15802
rect 14266 15750 14278 15802
rect 14330 15750 14342 15802
rect 14394 15750 14406 15802
rect 14458 15750 14470 15802
rect 14522 15750 14904 15802
rect 1104 15728 14904 15750
rect 934 15648 940 15700
rect 992 15688 998 15700
rect 1489 15691 1547 15697
rect 1489 15688 1501 15691
rect 992 15660 1501 15688
rect 992 15648 998 15660
rect 1489 15657 1501 15660
rect 1535 15657 1547 15691
rect 1489 15651 1547 15657
rect 7282 15648 7288 15700
rect 7340 15648 7346 15700
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 10468 15660 14289 15688
rect 10468 15648 10474 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 14 15444 20 15496
rect 72 15484 78 15496
rect 1949 15487 2007 15493
rect 1949 15484 1961 15487
rect 72 15456 1961 15484
rect 72 15444 78 15456
rect 1949 15453 1961 15456
rect 1995 15453 2007 15487
rect 1949 15447 2007 15453
rect 2682 15444 2688 15496
rect 2740 15444 2746 15496
rect 4614 15444 4620 15496
rect 4672 15444 4678 15496
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 9088 15456 9321 15484
rect 9088 15444 9094 15456
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11664 15456 11805 15484
rect 11664 15444 11670 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 13538 15444 13544 15496
rect 13596 15444 13602 15496
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15484 13967 15487
rect 15470 15484 15476 15496
rect 13955 15456 15476 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15416 1823 15419
rect 5718 15416 5724 15428
rect 1811 15388 5724 15416
rect 1811 15385 1823 15388
rect 1765 15379 1823 15385
rect 5718 15376 5724 15388
rect 5776 15376 5782 15428
rect 7561 15419 7619 15425
rect 7561 15385 7573 15419
rect 7607 15416 7619 15419
rect 7650 15416 7656 15428
rect 7607 15388 7656 15416
rect 7607 15385 7619 15388
rect 7561 15379 7619 15385
rect 7650 15376 7656 15388
rect 7708 15376 7714 15428
rect 13556 15416 13584 15444
rect 14185 15419 14243 15425
rect 14185 15416 14197 15419
rect 13556 15388 14197 15416
rect 14185 15385 14197 15388
rect 14231 15385 14243 15419
rect 14185 15379 14243 15385
rect 2130 15308 2136 15360
rect 2188 15308 2194 15360
rect 2866 15308 2872 15360
rect 2924 15308 2930 15360
rect 4798 15308 4804 15360
rect 4856 15308 4862 15360
rect 8754 15308 8760 15360
rect 8812 15348 8818 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8812 15320 9137 15348
rect 8812 15308 8818 15320
rect 9125 15317 9137 15320
rect 9171 15317 9183 15351
rect 9125 15311 9183 15317
rect 11882 15308 11888 15360
rect 11940 15308 11946 15360
rect 13722 15308 13728 15360
rect 13780 15308 13786 15360
rect 1104 15258 14904 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 14904 15258
rect 1104 15184 14904 15206
rect 14461 15147 14519 15153
rect 14461 15113 14473 15147
rect 14507 15144 14519 15147
rect 14826 15144 14832 15156
rect 14507 15116 14832 15144
rect 14507 15113 14519 15116
rect 14461 15107 14519 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13872 14980 14197 15008
rect 13872 14968 13878 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 1104 14714 14904 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 14214 14714
rect 14266 14662 14278 14714
rect 14330 14662 14342 14714
rect 14394 14662 14406 14714
rect 14458 14662 14470 14714
rect 14522 14662 14904 14714
rect 1104 14640 14904 14662
rect 1104 14170 14904 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 14904 14170
rect 1104 14096 14904 14118
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 7285 13923 7343 13929
rect 7285 13889 7297 13923
rect 7331 13920 7343 13923
rect 7926 13920 7932 13932
rect 7331 13892 7932 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 13964 13892 14197 13920
rect 13964 13880 13970 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 6546 13852 6552 13864
rect 1719 13824 6552 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 6546 13812 6552 13824
rect 6604 13812 6610 13864
rect 7374 13812 7380 13864
rect 7432 13812 7438 13864
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 14826 13852 14832 13864
rect 14507 13824 14832 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 14826 13812 14832 13824
rect 14884 13812 14890 13864
rect 7653 13787 7711 13793
rect 7653 13753 7665 13787
rect 7699 13784 7711 13787
rect 8202 13784 8208 13796
rect 7699 13756 8208 13784
rect 7699 13753 7711 13756
rect 7653 13747 7711 13753
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 9582 13716 9588 13728
rect 8536 13688 9588 13716
rect 8536 13676 8542 13688
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 1104 13626 14904 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 14214 13626
rect 14266 13574 14278 13626
rect 14330 13574 14342 13626
rect 14394 13574 14406 13626
rect 14458 13574 14470 13626
rect 14522 13574 14904 13626
rect 1104 13552 14904 13574
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 4798 13512 4804 13524
rect 4571 13484 4804 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 5442 13512 5448 13524
rect 5123 13484 5448 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 4816 13317 4844 13472
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 4264 13240 4292 13271
rect 5092 13240 5120 13475
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6546 13472 6552 13524
rect 6604 13512 6610 13524
rect 9490 13512 9496 13524
rect 6604 13484 9496 13512
rect 6604 13472 6610 13484
rect 9490 13472 9496 13484
rect 9548 13512 9554 13524
rect 9548 13484 10824 13512
rect 9548 13472 9554 13484
rect 8478 13444 8484 13456
rect 7484 13416 8484 13444
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5445 13379 5503 13385
rect 5445 13376 5457 13379
rect 5316 13348 5457 13376
rect 5316 13336 5322 13348
rect 5445 13345 5457 13348
rect 5491 13345 5503 13379
rect 5445 13339 5503 13345
rect 5905 13379 5963 13385
rect 5905 13345 5917 13379
rect 5951 13376 5963 13379
rect 5994 13376 6000 13388
rect 5951 13348 6000 13376
rect 5951 13345 5963 13348
rect 5905 13339 5963 13345
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 5350 13268 5356 13320
rect 5408 13308 5414 13320
rect 5537 13311 5595 13317
rect 5537 13308 5549 13311
rect 5408 13280 5549 13308
rect 5408 13268 5414 13280
rect 5537 13277 5549 13280
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 6546 13268 6552 13320
rect 6604 13268 6610 13320
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7484 13317 7512 13416
rect 8478 13404 8484 13416
rect 8536 13404 8542 13456
rect 9677 13447 9735 13453
rect 9677 13444 9689 13447
rect 8588 13416 9689 13444
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 8588 13385 8616 13416
rect 9677 13413 9689 13416
rect 9723 13413 9735 13447
rect 10410 13444 10416 13456
rect 9677 13407 9735 13413
rect 9968 13416 10416 13444
rect 8573 13379 8631 13385
rect 7800 13348 8524 13376
rect 7800 13336 7806 13348
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 6788 13280 7481 13308
rect 6788 13268 6794 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 8294 13268 8300 13320
rect 8352 13268 8358 13320
rect 8496 13317 8524 13348
rect 8573 13345 8585 13379
rect 8619 13345 8631 13379
rect 8573 13339 8631 13345
rect 9122 13336 9128 13388
rect 9180 13336 9186 13388
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 9968 13385 9996 13416
rect 10410 13404 10416 13416
rect 10468 13404 10474 13456
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9640 13348 9965 13376
rect 9640 13336 9646 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13376 10103 13379
rect 10091 13348 10548 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 9214 13308 9220 13320
rect 8527 13280 9220 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 4264 13212 5120 13240
rect 7926 13200 7932 13252
rect 7984 13240 7990 13252
rect 8021 13243 8079 13249
rect 8021 13240 8033 13243
rect 7984 13212 8033 13240
rect 7984 13200 7990 13212
rect 8021 13209 8033 13212
rect 8067 13240 8079 13243
rect 8404 13240 8432 13271
rect 9214 13268 9220 13280
rect 9272 13308 9278 13320
rect 9858 13308 9864 13320
rect 9272 13280 9864 13308
rect 9272 13268 9278 13280
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10410 13308 10416 13320
rect 10367 13280 10416 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 10520 13317 10548 13348
rect 10796 13317 10824 13484
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 10551 13280 10701 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 10042 13240 10048 13252
rect 8067 13212 8432 13240
rect 9600 13212 10048 13240
rect 8067 13209 8079 13212
rect 8021 13203 8079 13209
rect 4706 13132 4712 13184
rect 4764 13132 4770 13184
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 9600 13181 9628 13212
rect 10042 13200 10048 13212
rect 10100 13200 10106 13252
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 7892 13144 8125 13172
rect 7892 13132 7898 13144
rect 8113 13141 8125 13144
rect 8159 13141 8171 13175
rect 8113 13135 8171 13141
rect 9585 13175 9643 13181
rect 9585 13141 9597 13175
rect 9631 13141 9643 13175
rect 9585 13135 9643 13141
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9732 13144 10425 13172
rect 9732 13132 9738 13144
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 10413 13135 10471 13141
rect 1104 13082 14904 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 14904 13082
rect 1104 13008 14904 13030
rect 4706 12928 4712 12980
rect 4764 12928 4770 12980
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5215 12940 6914 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 4724 12900 4752 12928
rect 5077 12903 5135 12909
rect 5077 12900 5089 12903
rect 4356 12872 5089 12900
rect 4356 12841 4384 12872
rect 5077 12869 5089 12872
rect 5123 12869 5135 12903
rect 5077 12863 5135 12869
rect 5258 12860 5264 12912
rect 5316 12860 5322 12912
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 4448 12764 4476 12795
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 4764 12804 4997 12832
rect 4764 12792 4770 12804
rect 4985 12801 4997 12804
rect 5031 12832 5043 12835
rect 5350 12832 5356 12844
rect 5031 12804 5356 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 6886 12832 6914 12940
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 8018 12968 8024 12980
rect 7432 12940 8024 12968
rect 7432 12928 7438 12940
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 8294 12928 8300 12980
rect 8352 12928 8358 12980
rect 8842 12971 8900 12977
rect 8842 12937 8854 12971
rect 8888 12968 8900 12971
rect 9122 12968 9128 12980
rect 8888 12940 9128 12968
rect 8888 12937 8900 12940
rect 8842 12931 8900 12937
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9674 12928 9680 12980
rect 9732 12928 9738 12980
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10192 12940 10425 12968
rect 10192 12928 10198 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 8312 12900 8340 12928
rect 7484 12872 8340 12900
rect 8941 12903 8999 12909
rect 7484 12841 7512 12872
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6886 12804 7297 12832
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 4724 12764 4752 12792
rect 4448 12736 4752 12764
rect 7300 12764 7328 12795
rect 7668 12764 7696 12795
rect 7742 12792 7748 12844
rect 7800 12792 7806 12844
rect 7300 12736 7696 12764
rect 7852 12696 7880 12872
rect 8941 12869 8953 12903
rect 8987 12900 8999 12903
rect 9692 12900 9720 12928
rect 8987 12872 9720 12900
rect 8987 12869 8999 12872
rect 8941 12863 8999 12869
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 11517 12903 11575 12909
rect 11517 12900 11529 12903
rect 9916 12872 11529 12900
rect 9916 12860 9922 12872
rect 11517 12869 11529 12872
rect 11563 12869 11575 12903
rect 11517 12863 11575 12869
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8076 12804 8677 12832
rect 8076 12792 8082 12804
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 10962 12832 10968 12844
rect 10919 12804 10968 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 7944 12764 7972 12792
rect 8772 12764 8800 12795
rect 10962 12792 10968 12804
rect 11020 12832 11026 12844
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 11020 12804 12449 12832
rect 11020 12792 11026 12804
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12832 13415 12835
rect 13722 12832 13728 12844
rect 13403 12804 13728 12832
rect 13403 12801 13415 12804
rect 13357 12795 13415 12801
rect 7944 12736 8800 12764
rect 4816 12668 7880 12696
rect 8297 12699 8355 12705
rect 4816 12637 4844 12668
rect 8297 12665 8309 12699
rect 8343 12696 8355 12699
rect 8386 12696 8392 12708
rect 8343 12668 8392 12696
rect 8343 12665 8355 12668
rect 8297 12659 8355 12665
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 10597 12699 10655 12705
rect 10597 12665 10609 12699
rect 10643 12696 10655 12699
rect 11330 12696 11336 12708
rect 10643 12668 11336 12696
rect 10643 12665 10655 12668
rect 10597 12659 10655 12665
rect 11330 12656 11336 12668
rect 11388 12696 11394 12708
rect 13372 12696 13400 12795
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 11388 12668 13400 12696
rect 11388 12656 11394 12668
rect 4801 12631 4859 12637
rect 4801 12597 4813 12631
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 1104 12538 14904 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 14214 12538
rect 14266 12486 14278 12538
rect 14330 12486 14342 12538
rect 14394 12486 14406 12538
rect 14458 12486 14470 12538
rect 14522 12486 14904 12538
rect 1104 12464 14904 12486
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 5960 12260 9996 12288
rect 5960 12248 5966 12260
rect 9968 12232 9996 12260
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 6086 12180 6092 12232
rect 6144 12180 6150 12232
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 4724 12152 4752 12180
rect 6288 12152 6316 12183
rect 9950 12180 9956 12232
rect 10008 12180 10014 12232
rect 6362 12152 6368 12164
rect 4724 12124 6368 12152
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 13906 12152 13912 12164
rect 8812 12124 13912 12152
rect 8812 12112 8818 12124
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 6270 12044 6276 12096
rect 6328 12044 6334 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 11054 12084 11060 12096
rect 7248 12056 11060 12084
rect 7248 12044 7254 12056
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 1104 11994 14904 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 14904 11994
rect 1104 11920 14904 11942
rect 3878 11840 3884 11892
rect 3936 11880 3942 11892
rect 3936 11852 4568 11880
rect 3936 11840 3942 11852
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 4540 11812 4568 11852
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 4709 11883 4767 11889
rect 4709 11880 4721 11883
rect 4672 11852 4721 11880
rect 4672 11840 4678 11852
rect 4709 11849 4721 11852
rect 4755 11849 4767 11883
rect 4709 11843 4767 11849
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 6086 11880 6092 11892
rect 5583 11852 6092 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 8294 11880 8300 11892
rect 6196 11852 8300 11880
rect 5169 11815 5227 11821
rect 5169 11812 5181 11815
rect 1811 11784 4476 11812
rect 4540 11784 5181 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 3878 11704 3884 11756
rect 3936 11704 3942 11756
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4448 11676 4476 11784
rect 5169 11781 5181 11784
rect 5215 11781 5227 11815
rect 5169 11775 5227 11781
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 6196 11812 6224 11852
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 8754 11840 8760 11892
rect 8812 11840 8818 11892
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 10229 11883 10287 11889
rect 9539 11852 9904 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 5500 11784 6224 11812
rect 5500 11772 5506 11784
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11744 4675 11747
rect 4706 11744 4712 11756
rect 4663 11716 4712 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 4798 11704 4804 11756
rect 4856 11744 4862 11756
rect 5350 11744 5356 11756
rect 4856 11716 5356 11744
rect 4856 11704 4862 11716
rect 5350 11704 5356 11716
rect 5408 11704 5414 11756
rect 5552 11753 5580 11784
rect 6270 11772 6276 11824
rect 6328 11772 6334 11824
rect 7745 11815 7803 11821
rect 7745 11781 7757 11815
rect 7791 11812 7803 11815
rect 8772 11812 8800 11840
rect 9876 11821 9904 11852
rect 10229 11849 10241 11883
rect 10275 11880 10287 11883
rect 10275 11852 10640 11880
rect 10275 11849 10287 11852
rect 10229 11843 10287 11849
rect 7791 11784 8800 11812
rect 9861 11815 9919 11821
rect 7791 11781 7803 11784
rect 7745 11775 7803 11781
rect 9861 11781 9873 11815
rect 9907 11781 9919 11815
rect 9861 11775 9919 11781
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5736 11676 5764 11707
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 5994 11704 6000 11756
rect 6052 11704 6058 11756
rect 6288 11744 6316 11772
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 6288 11716 6653 11744
rect 6641 11713 6653 11716
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 7374 11744 7380 11756
rect 6779 11716 7380 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 6365 11679 6423 11685
rect 6365 11676 6377 11679
rect 4019 11648 4108 11676
rect 4448 11648 5672 11676
rect 5736 11648 6377 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 4080 11620 4108 11648
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 4801 11611 4859 11617
rect 4801 11608 4813 11611
rect 4120 11580 4813 11608
rect 4120 11568 4126 11580
rect 4801 11577 4813 11580
rect 4847 11577 4859 11611
rect 4801 11571 4859 11577
rect 5644 11540 5672 11648
rect 6365 11645 6377 11648
rect 6411 11645 6423 11679
rect 6365 11639 6423 11645
rect 6546 11636 6552 11688
rect 6604 11636 6610 11688
rect 6822 11636 6828 11688
rect 6880 11636 6886 11688
rect 6181 11611 6239 11617
rect 6181 11577 6193 11611
rect 6227 11608 6239 11611
rect 7760 11608 7788 11775
rect 9950 11772 9956 11824
rect 10008 11772 10014 11824
rect 10612 11821 10640 11852
rect 11054 11840 11060 11892
rect 11112 11840 11118 11892
rect 10597 11815 10655 11821
rect 10597 11781 10609 11815
rect 10643 11781 10655 11815
rect 10597 11775 10655 11781
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 6227 11580 7788 11608
rect 7852 11716 7941 11744
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 7190 11540 7196 11552
rect 5644 11512 7196 11540
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 7558 11500 7564 11552
rect 7616 11500 7622 11552
rect 7852 11540 7880 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8202 11704 8208 11756
rect 8260 11704 8266 11756
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11676 8079 11679
rect 8110 11676 8116 11688
rect 8067 11648 8116 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8312 11676 8340 11707
rect 9122 11704 9128 11756
rect 9180 11704 9186 11756
rect 9766 11753 9772 11756
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9733 11747 9772 11753
rect 9733 11713 9745 11747
rect 9733 11707 9772 11713
rect 8846 11676 8852 11688
rect 8312 11648 8852 11676
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 9140 11608 9168 11704
rect 9214 11636 9220 11688
rect 9272 11636 9278 11688
rect 9600 11676 9628 11707
rect 9766 11704 9772 11707
rect 9824 11704 9830 11756
rect 10042 11704 10048 11756
rect 10100 11753 10106 11756
rect 10100 11744 10108 11753
rect 10100 11716 10145 11744
rect 10100 11707 10108 11716
rect 10100 11704 10106 11707
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 11011 11716 11253 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11241 11713 11253 11716
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 9858 11676 9864 11688
rect 9600 11648 9864 11676
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 13814 11608 13820 11620
rect 7984 11580 9168 11608
rect 9508 11580 13820 11608
rect 7984 11568 7990 11580
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 7852 11512 8125 11540
rect 8113 11509 8125 11512
rect 8159 11540 8171 11543
rect 9508 11540 9536 11580
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 8159 11512 9536 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 1104 11450 14904 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 14214 11450
rect 14266 11398 14278 11450
rect 14330 11398 14342 11450
rect 14394 11398 14406 11450
rect 14458 11398 14470 11450
rect 14522 11398 14904 11450
rect 1104 11376 14904 11398
rect 5077 11339 5135 11345
rect 5077 11305 5089 11339
rect 5123 11336 5135 11339
rect 5626 11336 5632 11348
rect 5123 11308 5632 11336
rect 5123 11305 5135 11308
rect 5077 11299 5135 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6086 11296 6092 11348
rect 6144 11296 6150 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6546 11336 6552 11348
rect 6503 11308 6552 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6546 11296 6552 11308
rect 6604 11336 6610 11348
rect 7282 11336 7288 11348
rect 6604 11308 7288 11336
rect 6604 11296 6610 11308
rect 7282 11296 7288 11308
rect 7340 11336 7346 11348
rect 7340 11308 8248 11336
rect 7340 11296 7346 11308
rect 4080 11240 5396 11268
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4080 11132 4108 11240
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 4212 11172 4629 11200
rect 4212 11160 4218 11172
rect 4617 11169 4629 11172
rect 4663 11200 4675 11203
rect 4663 11172 5212 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 3936 11104 4537 11132
rect 3936 11092 3942 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 5184 11141 5212 11172
rect 5368 11141 5396 11240
rect 6104 11141 6132 11296
rect 7208 11240 8156 11268
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 7208 11132 7236 11240
rect 6089 11095 6147 11101
rect 6196 11104 7236 11132
rect 4908 11064 4936 11095
rect 5261 11067 5319 11073
rect 4908 11036 5212 11064
rect 5184 10996 5212 11036
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 6196 11064 6224 11104
rect 5307 11036 6224 11064
rect 6273 11067 6331 11073
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 6273 11033 6285 11067
rect 6319 11064 6331 11067
rect 6362 11064 6368 11076
rect 6319 11036 6368 11064
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 7208 11064 7236 11104
rect 7282 11092 7288 11144
rect 7340 11092 7346 11144
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7834 11132 7840 11144
rect 7607 11104 7840 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8128 11141 8156 11240
rect 8220 11144 8248 11308
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 9769 11339 9827 11345
rect 9769 11336 9781 11339
rect 9272 11308 9781 11336
rect 9272 11296 9278 11308
rect 9769 11305 9781 11308
rect 9815 11305 9827 11339
rect 9769 11299 9827 11305
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10836 11308 10885 11336
rect 10836 11296 10842 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 10873 11299 10931 11305
rect 11330 11296 11336 11348
rect 11388 11296 11394 11348
rect 8389 11271 8447 11277
rect 8389 11237 8401 11271
rect 8435 11268 8447 11271
rect 9674 11268 9680 11280
rect 8435 11240 9680 11268
rect 8435 11237 8447 11240
rect 8389 11231 8447 11237
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 8352 11172 14289 11200
rect 8352 11160 8358 11172
rect 14277 11169 14289 11172
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 8076 11104 8125 11132
rect 8076 11092 8082 11104
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 8202 11092 8208 11144
rect 8260 11092 8266 11144
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10594 11132 10600 11144
rect 9640 11104 10600 11132
rect 9640 11092 9646 11104
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 7377 11067 7435 11073
rect 7377 11064 7389 11067
rect 7208 11036 7389 11064
rect 7377 11033 7389 11036
rect 7423 11033 7435 11067
rect 7377 11027 7435 11033
rect 7745 11067 7803 11073
rect 7745 11033 7757 11067
rect 7791 11064 7803 11067
rect 8570 11064 8576 11076
rect 7791 11036 8576 11064
rect 7791 11033 7803 11036
rect 7745 11027 7803 11033
rect 8570 11024 8576 11036
rect 8628 11064 8634 11076
rect 9125 11067 9183 11073
rect 9125 11064 9137 11067
rect 8628 11036 9137 11064
rect 8628 11024 8634 11036
rect 9125 11033 9137 11036
rect 9171 11033 9183 11067
rect 11072 11064 11100 11095
rect 11146 11092 11152 11144
rect 11204 11092 11210 11144
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11422 11132 11428 11144
rect 11296 11104 11428 11132
rect 11296 11092 11302 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 14599 11104 14964 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 14936 11076 14964 11104
rect 11698 11064 11704 11076
rect 9125 11027 9183 11033
rect 9232 11036 11704 11064
rect 6546 10996 6552 11008
rect 5184 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10996 6610 11008
rect 9232 10996 9260 11036
rect 11698 11024 11704 11036
rect 11756 11024 11762 11076
rect 14918 11024 14924 11076
rect 14976 11024 14982 11076
rect 6604 10968 9260 10996
rect 6604 10956 6610 10968
rect 1104 10906 14904 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 14904 10906
rect 1104 10832 14904 10854
rect 4617 10795 4675 10801
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 4798 10792 4804 10804
rect 4663 10764 4804 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 8047 10795 8105 10801
rect 8047 10761 8059 10795
rect 8093 10792 8105 10795
rect 8202 10792 8208 10804
rect 8093 10764 8208 10792
rect 8093 10761 8105 10764
rect 8047 10755 8105 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 11146 10752 11152 10804
rect 11204 10752 11210 10804
rect 7282 10684 7288 10736
rect 7340 10724 7346 10736
rect 7834 10724 7840 10736
rect 7340 10696 7840 10724
rect 7340 10684 7346 10696
rect 7834 10684 7840 10696
rect 7892 10684 7898 10736
rect 4154 10656 4160 10668
rect 2240 10628 4160 10656
rect 2240 10532 2268 10628
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4387 10628 4537 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4525 10625 4537 10628
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 6914 10656 6920 10668
rect 4755 10628 6920 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3936 10560 3985 10588
rect 3936 10548 3942 10560
rect 3973 10557 3985 10560
rect 4019 10557 4031 10591
rect 3973 10551 4031 10557
rect 2222 10480 2228 10532
rect 2280 10480 2286 10532
rect 4540 10520 4568 10619
rect 6914 10616 6920 10628
rect 6972 10656 6978 10668
rect 6972 10628 9674 10656
rect 6972 10616 6978 10628
rect 9646 10588 9674 10628
rect 10962 10616 10968 10668
rect 11020 10656 11026 10668
rect 11057 10659 11115 10665
rect 11057 10656 11069 10659
rect 11020 10628 11069 10656
rect 11020 10616 11026 10628
rect 11057 10625 11069 10628
rect 11103 10625 11115 10659
rect 11057 10619 11115 10625
rect 11241 10659 11299 10665
rect 11241 10625 11253 10659
rect 11287 10656 11299 10659
rect 11606 10656 11612 10668
rect 11287 10628 11612 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11256 10588 11284 10619
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 9646 10560 11284 10588
rect 4798 10520 4804 10532
rect 4540 10492 4804 10520
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 9306 10520 9312 10532
rect 6288 10492 9312 10520
rect 6288 10464 6316 10492
rect 9306 10480 9312 10492
rect 9364 10480 9370 10532
rect 6270 10412 6276 10464
rect 6328 10412 6334 10464
rect 8018 10412 8024 10464
rect 8076 10412 8082 10464
rect 8205 10455 8263 10461
rect 8205 10421 8217 10455
rect 8251 10452 8263 10455
rect 8294 10452 8300 10464
rect 8251 10424 8300 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 1104 10362 14904 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 14214 10362
rect 14266 10310 14278 10362
rect 14330 10310 14342 10362
rect 14394 10310 14406 10362
rect 14458 10310 14470 10362
rect 14522 10310 14904 10362
rect 1104 10288 14904 10310
rect 8294 10208 8300 10260
rect 8352 10208 8358 10260
rect 8478 10208 8484 10260
rect 8536 10208 8542 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9548 10220 9674 10248
rect 9548 10208 9554 10220
rect 5442 10180 5448 10192
rect 4356 10152 5448 10180
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4213 10047 4271 10053
rect 4213 10013 4225 10047
rect 4259 10044 4271 10047
rect 4356 10044 4384 10152
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 6273 10183 6331 10189
rect 6273 10149 6285 10183
rect 6319 10180 6331 10183
rect 7466 10180 7472 10192
rect 6319 10152 7472 10180
rect 6319 10149 6331 10152
rect 6273 10143 6331 10149
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 4798 10112 4804 10124
rect 4448 10084 4804 10112
rect 4448 10053 4476 10084
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 5644 10084 6377 10112
rect 4259 10016 4384 10044
rect 4433 10047 4491 10053
rect 4259 10013 4271 10016
rect 4213 10007 4271 10013
rect 4433 10013 4445 10047
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4571 10047 4629 10053
rect 4571 10013 4583 10047
rect 4617 10044 4629 10047
rect 5258 10044 5264 10056
rect 4617 10016 5264 10044
rect 4617 10013 4629 10016
rect 4571 10007 4629 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5644 10053 5672 10084
rect 6365 10081 6377 10084
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6472 10084 6684 10112
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5722 10047 5780 10053
rect 5722 10013 5734 10047
rect 5768 10013 5780 10047
rect 5722 10007 5780 10013
rect 4338 9936 4344 9988
rect 4396 9936 4402 9988
rect 5736 9976 5764 10007
rect 6086 10004 6092 10056
rect 6144 10053 6150 10056
rect 6144 10047 6193 10053
rect 6144 10013 6147 10047
rect 6181 10044 6193 10047
rect 6472 10044 6500 10084
rect 6656 10056 6684 10084
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 8312 10121 8340 10208
rect 9646 10180 9674 10220
rect 9858 10208 9864 10260
rect 9916 10208 9922 10260
rect 10134 10208 10140 10260
rect 10192 10208 10198 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10962 10248 10968 10260
rect 10284 10220 10968 10248
rect 10284 10208 10290 10220
rect 10962 10208 10968 10220
rect 11020 10248 11026 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 11020 10220 11069 10248
rect 11020 10208 11026 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 9380 10152 10824 10180
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 8297 10115 8355 10121
rect 6871 10084 8156 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 6181 10016 6500 10044
rect 6181 10013 6193 10016
rect 6144 10007 6193 10013
rect 6144 10004 6150 10007
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 4632 9948 5764 9976
rect 4632 9920 4660 9948
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 5905 9979 5963 9985
rect 5905 9976 5917 9979
rect 5868 9948 5917 9976
rect 5868 9936 5874 9948
rect 5905 9945 5917 9948
rect 5951 9945 5963 9979
rect 5905 9939 5963 9945
rect 5997 9979 6055 9985
rect 5997 9945 6009 9979
rect 6043 9976 6055 9979
rect 6270 9976 6276 9988
rect 6043 9948 6276 9976
rect 6043 9945 6055 9948
rect 5997 9939 6055 9945
rect 6270 9936 6276 9948
rect 6328 9936 6334 9988
rect 6362 9936 6368 9988
rect 6420 9976 6426 9988
rect 6840 9976 6868 10075
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 7181 10047 7239 10053
rect 7181 10044 7193 10047
rect 7116 10016 7193 10044
rect 6420 9948 6868 9976
rect 6932 9976 6960 10004
rect 7116 9976 7144 10016
rect 7181 10013 7193 10016
rect 7227 10013 7239 10047
rect 7181 10007 7239 10013
rect 7282 10004 7288 10056
rect 7340 10004 7346 10056
rect 7576 10053 7604 10084
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 7561 10047 7619 10053
rect 7423 10016 7512 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 6932 9948 7144 9976
rect 7484 9976 7512 10016
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 8128 10044 8156 10084
rect 8297 10081 8309 10115
rect 8343 10081 8355 10115
rect 9380 10112 9408 10152
rect 8297 10075 8355 10081
rect 8404 10084 9408 10112
rect 8404 10044 8432 10084
rect 8128 10016 8432 10044
rect 7561 10007 7619 10013
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 9214 10004 9220 10056
rect 9272 10004 9278 10056
rect 9380 10053 9408 10084
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 9640 10084 10456 10112
rect 9640 10072 9646 10084
rect 9365 10047 9423 10053
rect 9365 10013 9377 10047
rect 9411 10013 9423 10047
rect 9365 10007 9423 10013
rect 9723 10047 9781 10053
rect 9723 10013 9735 10047
rect 9769 10044 9781 10047
rect 9858 10044 9864 10056
rect 9769 10016 9864 10044
rect 9769 10013 9781 10016
rect 9723 10007 9781 10013
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10428 10053 10456 10084
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 7926 9976 7932 9988
rect 7484 9948 7932 9976
rect 6420 9936 6426 9948
rect 7926 9936 7932 9948
rect 7984 9936 7990 9988
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 9493 9979 9551 9985
rect 9493 9976 9505 9979
rect 8812 9948 9505 9976
rect 8812 9936 8818 9948
rect 9493 9945 9505 9948
rect 9539 9945 9551 9979
rect 9493 9939 9551 9945
rect 9585 9979 9643 9985
rect 9585 9945 9597 9979
rect 9631 9976 9643 9979
rect 10226 9976 10232 9988
rect 9631 9948 10232 9976
rect 9631 9945 9643 9948
rect 9585 9939 9643 9945
rect 4614 9868 4620 9920
rect 4672 9868 4678 9920
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 6822 9908 6828 9920
rect 4755 9880 6828 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 8018 9868 8024 9920
rect 8076 9868 8082 9920
rect 9508 9908 9536 9939
rect 10226 9936 10232 9948
rect 10284 9936 10290 9988
rect 10042 9908 10048 9920
rect 9508 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 10428 9908 10456 10007
rect 10520 9976 10548 10007
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 10796 10053 10824 10152
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10044 11299 10047
rect 11330 10044 11336 10056
rect 11287 10016 11336 10044
rect 11287 10013 11299 10016
rect 11241 10007 11299 10013
rect 11256 9976 11284 10007
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 11440 9976 11468 10004
rect 11974 9976 11980 9988
rect 10520 9948 11284 9976
rect 11348 9948 11980 9976
rect 11348 9908 11376 9948
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 10428 9880 11376 9908
rect 1104 9818 14904 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 14904 9818
rect 1104 9744 14904 9766
rect 3697 9707 3755 9713
rect 3697 9673 3709 9707
rect 3743 9704 3755 9707
rect 4062 9704 4068 9716
rect 3743 9676 4068 9704
rect 3743 9673 3755 9676
rect 3697 9667 3755 9673
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 5810 9704 5816 9716
rect 4396 9676 5816 9704
rect 4396 9664 4402 9676
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 6730 9704 6736 9716
rect 6656 9676 6736 9704
rect 4249 9639 4307 9645
rect 4249 9605 4261 9639
rect 4295 9636 4307 9639
rect 6362 9636 6368 9648
rect 4295 9608 6368 9636
rect 4295 9605 4307 9608
rect 4249 9599 4307 9605
rect 6362 9596 6368 9608
rect 6420 9636 6426 9648
rect 6656 9645 6684 9676
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 7837 9707 7895 9713
rect 7837 9673 7849 9707
rect 7883 9704 7895 9707
rect 8018 9704 8024 9716
rect 7883 9676 8024 9704
rect 7883 9673 7895 9676
rect 7837 9667 7895 9673
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 9214 9664 9220 9716
rect 9272 9664 9278 9716
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 10137 9707 10195 9713
rect 10137 9704 10149 9707
rect 9640 9676 10149 9704
rect 9640 9664 9646 9676
rect 10137 9673 10149 9676
rect 10183 9673 10195 9707
rect 10137 9667 10195 9673
rect 6641 9639 6699 9645
rect 6420 9608 6592 9636
rect 6420 9596 6426 9608
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3804 9540 3985 9568
rect 3804 9432 3832 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 4706 9568 4712 9580
rect 4387 9540 4712 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 4706 9528 4712 9540
rect 4764 9568 4770 9580
rect 6086 9568 6092 9580
rect 4764 9540 6092 9568
rect 4764 9528 4770 9540
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9537 6515 9571
rect 6564 9568 6592 9608
rect 6641 9605 6653 9639
rect 6687 9605 6699 9639
rect 6641 9599 6699 9605
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 6880 9608 9628 9636
rect 6880 9596 6886 9608
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 6564 9540 6745 9568
rect 6457 9531 6515 9537
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6840 9540 7420 9568
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 4614 9500 4620 9512
rect 3936 9472 4620 9500
rect 3936 9460 3942 9472
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 6472 9500 6500 9531
rect 6840 9500 6868 9540
rect 5224 9472 6868 9500
rect 5224 9460 5230 9472
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 7392 9500 7420 9540
rect 7466 9528 7472 9580
rect 7524 9528 7530 9580
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 9490 9568 9496 9580
rect 7984 9540 9496 9568
rect 7984 9528 7990 9540
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9600 9568 9628 9608
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 9950 9636 9956 9648
rect 9732 9608 9956 9636
rect 9732 9596 9738 9608
rect 9950 9596 9956 9608
rect 10008 9596 10014 9648
rect 10226 9634 10232 9686
rect 10284 9674 10290 9686
rect 10284 9646 10364 9674
rect 10284 9634 10290 9646
rect 9600 9540 9904 9568
rect 7392 9472 8248 9500
rect 6733 9435 6791 9441
rect 3804 9404 4844 9432
rect 4816 9376 4844 9404
rect 6733 9401 6745 9435
rect 6779 9432 6791 9435
rect 7024 9432 7052 9460
rect 6779 9404 7052 9432
rect 8021 9435 8079 9441
rect 6779 9401 6791 9404
rect 6733 9395 6791 9401
rect 8021 9401 8033 9435
rect 8067 9432 8079 9435
rect 8110 9432 8116 9444
rect 8067 9404 8116 9432
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 8220 9376 8248 9472
rect 9306 9460 9312 9512
rect 9364 9500 9370 9512
rect 9876 9509 9904 9540
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 10100 9540 10149 9568
rect 10100 9528 10106 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 10336 9577 10364 9646
rect 10428 9608 11100 9636
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9364 9472 9413 9500
rect 9364 9460 9370 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10428 9500 10456 9608
rect 11072 9580 11100 9608
rect 10505 9571 10563 9577
rect 10505 9537 10517 9571
rect 10551 9568 10563 9571
rect 10962 9568 10968 9580
rect 10551 9540 10968 9568
rect 10551 9537 10563 9540
rect 10505 9531 10563 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11054 9528 11060 9580
rect 11112 9528 11118 9580
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11698 9568 11704 9580
rect 11296 9540 11704 9568
rect 11296 9528 11302 9540
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 11882 9528 11888 9580
rect 11940 9528 11946 9580
rect 9907 9472 10456 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 9784 9432 9812 9463
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 11977 9503 12035 9509
rect 11977 9500 11989 9503
rect 10836 9472 11989 9500
rect 10836 9460 10842 9472
rect 11977 9469 11989 9472
rect 12023 9500 12035 9503
rect 12802 9500 12808 9512
rect 12023 9472 12808 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 10796 9432 10824 9460
rect 9784 9404 10824 9432
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 4338 9364 4344 9376
rect 3752 9336 4344 9364
rect 3752 9324 3758 9336
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4798 9324 4804 9376
rect 4856 9324 4862 9376
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7800 9336 7849 9364
rect 7800 9324 7806 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8202 9324 8208 9376
rect 8260 9324 8266 9376
rect 10318 9324 10324 9376
rect 10376 9324 10382 9376
rect 11514 9324 11520 9376
rect 11572 9324 11578 9376
rect 1104 9274 14904 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 14214 9274
rect 14266 9222 14278 9274
rect 14330 9222 14342 9274
rect 14394 9222 14406 9274
rect 14458 9222 14470 9274
rect 14522 9222 14904 9274
rect 1104 9200 14904 9222
rect 6914 9160 6920 9172
rect 2746 9132 6920 9160
rect 2746 9024 2774 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7650 9120 7656 9172
rect 7708 9169 7714 9172
rect 7708 9163 7757 9169
rect 7708 9129 7711 9163
rect 7745 9129 7757 9163
rect 7708 9123 7757 9129
rect 7708 9120 7714 9123
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10226 9160 10232 9172
rect 10100 9132 10232 9160
rect 10100 9120 10106 9132
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 10778 9120 10784 9172
rect 10836 9120 10842 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 10928 9132 11192 9160
rect 10928 9120 10934 9132
rect 4338 9092 4344 9104
rect 3988 9064 4344 9092
rect 3988 9033 4016 9064
rect 4338 9052 4344 9064
rect 4396 9092 4402 9104
rect 4396 9064 5488 9092
rect 4396 9052 4402 9064
rect 1780 8996 2774 9024
rect 3973 9027 4031 9033
rect 1780 8965 1808 8996
rect 3973 8993 3985 9027
rect 4019 8993 4031 9027
rect 5350 9024 5356 9036
rect 3973 8987 4031 8993
rect 4172 8996 5356 9024
rect 4172 8965 4200 8996
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5460 8968 5488 9064
rect 5718 9052 5724 9104
rect 5776 9092 5782 9104
rect 6822 9092 6828 9104
rect 5776 9064 6828 9092
rect 5776 9052 5782 9064
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 7208 9092 7236 9120
rect 7837 9095 7895 9101
rect 7837 9092 7849 9095
rect 7208 9064 7849 9092
rect 7837 9061 7849 9064
rect 7883 9061 7895 9095
rect 7837 9055 7895 9061
rect 8202 9052 8208 9104
rect 8260 9092 8266 9104
rect 8260 9064 9812 9092
rect 8260 9052 8266 9064
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 6748 8996 7941 9024
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 4614 8965 4620 8968
rect 4581 8959 4620 8965
rect 4581 8925 4593 8959
rect 4581 8919 4620 8925
rect 4614 8916 4620 8919
rect 4672 8916 4678 8968
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 4939 8959 4997 8965
rect 4939 8925 4951 8959
rect 4985 8956 4997 8959
rect 5166 8956 5172 8968
rect 4985 8928 5172 8956
rect 4985 8925 4997 8928
rect 4939 8919 4997 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 5442 8956 5448 8968
rect 5307 8928 5448 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 6546 8956 6552 8968
rect 5684 8928 6552 8956
rect 5684 8916 5690 8928
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 4801 8891 4859 8897
rect 4801 8888 4813 8891
rect 1397 8851 1455 8857
rect 4356 8860 4813 8888
rect 4356 8829 4384 8860
rect 4801 8857 4813 8860
rect 4847 8888 4859 8891
rect 5350 8888 5356 8900
rect 4847 8860 5356 8888
rect 4847 8857 4859 8860
rect 4801 8851 4859 8857
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 6656 8832 6684 8919
rect 6748 8832 6776 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 7558 8916 7564 8968
rect 7616 8916 7622 8968
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8343 8928 9045 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 6840 8888 6868 8916
rect 9416 8888 9444 8919
rect 6840 8860 9444 8888
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8789 4399 8823
rect 4341 8783 4399 8789
rect 5077 8823 5135 8829
rect 5077 8789 5089 8823
rect 5123 8820 5135 8823
rect 5442 8820 5448 8832
rect 5123 8792 5448 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 5810 8780 5816 8832
rect 5868 8780 5874 8832
rect 6638 8780 6644 8832
rect 6696 8780 6702 8832
rect 6730 8780 6736 8832
rect 6788 8780 6794 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7742 8820 7748 8832
rect 6972 8792 7748 8820
rect 6972 8780 6978 8792
rect 7742 8780 7748 8792
rect 7800 8820 7806 8832
rect 9692 8820 9720 8919
rect 9784 8900 9812 9064
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9916 8928 10149 8956
rect 9916 8916 9922 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 9766 8848 9772 8900
rect 9824 8888 9830 8900
rect 10689 8891 10747 8897
rect 9824 8860 10456 8888
rect 9824 8848 9830 8860
rect 7800 8792 9720 8820
rect 7800 8780 7806 8792
rect 10318 8780 10324 8832
rect 10376 8780 10382 8832
rect 10428 8820 10456 8860
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 10796 8888 10824 9120
rect 11057 9095 11115 9101
rect 11057 9061 11069 9095
rect 11103 9061 11115 9095
rect 11057 9055 11115 9061
rect 11072 8956 11100 9055
rect 11164 9024 11192 9132
rect 11514 9120 11520 9172
rect 11572 9120 11578 9172
rect 11882 9024 11888 9036
rect 11164 8996 11888 9024
rect 11882 8984 11888 8996
rect 11940 9024 11946 9036
rect 11940 8996 13216 9024
rect 11940 8984 11946 8996
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10919 8925 10977 8931
rect 11072 8928 11345 8956
rect 10919 8922 10931 8925
rect 10735 8860 10824 8888
rect 10904 8891 10931 8922
rect 10965 8891 10977 8925
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11514 8916 11520 8968
rect 11572 8916 11578 8968
rect 12802 8916 12808 8968
rect 12860 8916 12866 8968
rect 13188 8965 13216 8996
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13262 8956 13268 8968
rect 13219 8928 13268 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 10904 8888 10977 8891
rect 10904 8860 11008 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 10980 8832 11008 8860
rect 11790 8848 11796 8900
rect 11848 8848 11854 8900
rect 10962 8820 10968 8832
rect 10428 8792 10968 8820
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 12158 8780 12164 8832
rect 12216 8780 12222 8832
rect 1104 8730 14904 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 14904 8730
rect 1104 8656 14904 8678
rect 4062 8576 4068 8628
rect 4120 8576 4126 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4430 8616 4436 8628
rect 4203 8588 4436 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 5261 8619 5319 8625
rect 4939 8588 5120 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 3513 8551 3571 8557
rect 3513 8517 3525 8551
rect 3559 8548 3571 8551
rect 3786 8548 3792 8560
rect 3559 8520 3792 8548
rect 3559 8517 3571 8520
rect 3513 8511 3571 8517
rect 3786 8508 3792 8520
rect 3844 8548 3850 8560
rect 4080 8548 4108 8576
rect 4338 8548 4344 8560
rect 3844 8520 4108 8548
rect 4172 8520 4344 8548
rect 3844 8508 3850 8520
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4172 8480 4200 8520
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 4111 8452 4200 8480
rect 4249 8483 4307 8489
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 4798 8480 4804 8492
rect 4295 8452 4804 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5000 8412 5028 8443
rect 3436 8384 5028 8412
rect 3436 8288 3464 8384
rect 5092 8344 5120 8588
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 5534 8616 5540 8628
rect 5307 8588 5540 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5810 8576 5816 8628
rect 5868 8576 5874 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 7374 8576 7380 8628
rect 7432 8616 7438 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 7432 8588 7481 8616
rect 7432 8576 7438 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 7469 8579 7527 8585
rect 5350 8508 5356 8560
rect 5408 8508 5414 8560
rect 5442 8508 5448 8560
rect 5500 8508 5506 8560
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5368 8480 5396 8508
rect 5215 8452 5396 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5460 8412 5488 8508
rect 5828 8480 5856 8576
rect 6546 8508 6552 8560
rect 6604 8548 6610 8560
rect 7484 8548 7512 8579
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 7708 8588 8953 8616
rect 7708 8576 7714 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 9582 8616 9588 8628
rect 8941 8579 8999 8585
rect 9232 8588 9588 8616
rect 9232 8557 9260 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 11146 8616 11152 8628
rect 10336 8588 11152 8616
rect 9217 8551 9275 8557
rect 6604 8520 7420 8548
rect 7484 8520 7696 8548
rect 6604 8508 6610 8520
rect 6825 8483 6883 8489
rect 6825 8480 6837 8483
rect 5828 8452 6837 8480
rect 6825 8449 6837 8452
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 7098 8440 7104 8492
rect 7156 8440 7162 8492
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 5460 8384 7021 8412
rect 7009 8381 7021 8384
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7190 8372 7196 8424
rect 7248 8372 7254 8424
rect 7392 8421 7420 8520
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7668 8489 7696 8520
rect 9217 8517 9229 8551
rect 9263 8517 9275 8551
rect 10336 8548 10364 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 11790 8616 11796 8628
rect 11563 8588 11796 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 11940 8588 13952 8616
rect 11940 8576 11946 8588
rect 12158 8548 12164 8560
rect 9217 8511 9275 8517
rect 9600 8520 10364 8548
rect 10704 8520 12164 8548
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7524 8452 7573 8480
rect 7524 8440 7530 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 9122 8440 9128 8492
rect 9180 8440 9186 8492
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8381 7435 8415
rect 9324 8412 9352 8443
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9600 8489 9628 8520
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9456 8452 9505 8480
rect 9456 8440 9462 8452
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 9766 8440 9772 8492
rect 9824 8440 9830 8492
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 10008 8452 10149 8480
rect 10008 8440 10014 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10515 8489 10573 8495
rect 10704 8492 10732 8520
rect 10413 8483 10471 8489
rect 10413 8480 10425 8483
rect 10336 8452 10425 8480
rect 9674 8412 9680 8424
rect 9324 8384 9680 8412
rect 7377 8375 7435 8381
rect 9508 8356 9536 8384
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9784 8412 9812 8440
rect 10244 8412 10272 8440
rect 9784 8384 10272 8412
rect 6546 8344 6552 8356
rect 4172 8316 6552 8344
rect 3418 8236 3424 8288
rect 3476 8236 3482 8288
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4172 8276 4200 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 6840 8316 7297 8344
rect 6840 8288 6868 8316
rect 7285 8313 7297 8316
rect 7331 8313 7343 8347
rect 7285 8307 7343 8313
rect 7837 8347 7895 8353
rect 7837 8313 7849 8347
rect 7883 8344 7895 8347
rect 9490 8344 9496 8356
rect 7883 8316 9496 8344
rect 7883 8313 7895 8316
rect 7837 8307 7895 8313
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 9950 8304 9956 8356
rect 10008 8304 10014 8356
rect 10336 8344 10364 8452
rect 10413 8449 10425 8452
rect 10459 8449 10471 8483
rect 10515 8455 10527 8489
rect 10561 8486 10573 8489
rect 10561 8480 10640 8486
rect 10686 8480 10692 8492
rect 10561 8458 10692 8480
rect 10561 8455 10573 8458
rect 10515 8449 10573 8455
rect 10612 8452 10692 8458
rect 10413 8443 10471 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 11808 8489 11836 8520
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 12802 8480 12808 8492
rect 12115 8452 12808 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13924 8489 13952 8588
rect 14458 8508 14464 8560
rect 14516 8508 14522 8560
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 10336 8316 10640 8344
rect 3936 8248 4200 8276
rect 5077 8279 5135 8285
rect 3936 8236 3942 8248
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5166 8276 5172 8288
rect 5123 8248 5172 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 6822 8276 6828 8288
rect 5316 8248 6828 8276
rect 5316 8236 5322 8248
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 10612 8276 10640 8316
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11238 8344 11244 8356
rect 10744 8316 11244 8344
rect 10744 8304 10750 8316
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 11606 8344 11612 8356
rect 11388 8316 11612 8344
rect 11388 8304 11394 8316
rect 11606 8304 11612 8316
rect 11664 8344 11670 8356
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 11664 8316 11989 8344
rect 11664 8304 11670 8316
rect 11977 8313 11989 8316
rect 12023 8313 12035 8347
rect 11977 8307 12035 8313
rect 10962 8276 10968 8288
rect 10612 8248 10968 8276
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 1104 8186 14904 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 14214 8186
rect 14266 8134 14278 8186
rect 14330 8134 14342 8186
rect 14394 8134 14406 8186
rect 14458 8134 14470 8186
rect 14522 8134 14904 8186
rect 1104 8112 14904 8134
rect 6546 8032 6552 8084
rect 6604 8032 6610 8084
rect 8386 8032 8392 8084
rect 8444 8032 8450 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9180 8044 9413 8072
rect 9180 8032 9186 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 8004 4399 8007
rect 5166 8004 5172 8016
rect 4387 7976 5172 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 4433 7939 4491 7945
rect 3476 7908 4016 7936
rect 3476 7896 3482 7908
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 2961 7871 3019 7877
rect 2961 7868 2973 7871
rect 2924 7840 2973 7868
rect 2924 7828 2930 7840
rect 2961 7837 2973 7840
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3878 7828 3884 7880
rect 3936 7828 3942 7880
rect 3988 7877 4016 7908
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 5258 7936 5264 7948
rect 4479 7908 5264 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 7466 7936 7472 7948
rect 6472 7908 7472 7936
rect 6472 7880 6500 7908
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7892 7908 8125 7936
rect 7892 7896 7898 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 8202 7896 8208 7948
rect 8260 7896 8266 7948
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7936 8355 7939
rect 8404 7936 8432 8032
rect 8754 7936 8760 7948
rect 8343 7908 8760 7936
rect 8343 7905 8355 7908
rect 8297 7899 8355 7905
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 10502 7936 10508 7948
rect 9600 7908 10508 7936
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4062 7868 4068 7880
rect 4019 7840 4068 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 6822 7868 6828 7880
rect 6687 7840 6828 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7190 7868 7196 7880
rect 7055 7840 7196 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 2777 7803 2835 7809
rect 2777 7769 2789 7803
rect 2823 7800 2835 7803
rect 3896 7800 3924 7828
rect 2823 7772 3924 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 5368 7800 5396 7828
rect 7024 7800 7052 7831
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 7852 7840 8401 7868
rect 4488 7772 5396 7800
rect 6656 7772 7052 7800
rect 4488 7760 4494 7772
rect 6656 7744 6684 7772
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 4614 7732 4620 7744
rect 3568 7704 4620 7732
rect 3568 7692 3574 7704
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 4798 7732 4804 7744
rect 4755 7704 4804 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 4798 7692 4804 7704
rect 4856 7732 4862 7744
rect 5350 7732 5356 7744
rect 4856 7704 5356 7732
rect 4856 7692 4862 7704
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 6638 7692 6644 7744
rect 6696 7692 6702 7744
rect 6825 7735 6883 7741
rect 6825 7701 6837 7735
rect 6871 7732 6883 7735
rect 6914 7732 6920 7744
rect 6871 7704 6920 7732
rect 6871 7701 6883 7704
rect 6825 7695 6883 7701
rect 6914 7692 6920 7704
rect 6972 7732 6978 7744
rect 7852 7732 7880 7840
rect 8389 7837 8401 7840
rect 8435 7868 8447 7871
rect 8846 7868 8852 7880
rect 8435 7840 8852 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 8846 7828 8852 7840
rect 8904 7868 8910 7880
rect 9306 7868 9312 7880
rect 8904 7840 9312 7868
rect 8904 7828 8910 7840
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9600 7877 9628 7908
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 12860 7908 13093 7936
rect 12860 7896 12866 7908
rect 13081 7905 13093 7908
rect 13127 7905 13139 7939
rect 13081 7899 13139 7905
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10042 7868 10048 7880
rect 9907 7840 10048 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 12253 7803 12311 7809
rect 12253 7800 12265 7803
rect 9646 7772 12265 7800
rect 6972 7704 7880 7732
rect 6972 7692 6978 7704
rect 7926 7692 7932 7744
rect 7984 7692 7990 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 9030 7732 9036 7744
rect 8260 7704 9036 7732
rect 8260 7692 8266 7704
rect 9030 7692 9036 7704
rect 9088 7732 9094 7744
rect 9646 7732 9674 7772
rect 12253 7769 12265 7772
rect 12299 7769 12311 7803
rect 13188 7800 13216 7854
rect 13188 7772 13308 7800
rect 12253 7763 12311 7769
rect 13280 7744 13308 7772
rect 9088 7704 9674 7732
rect 9088 7692 9094 7704
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 11790 7732 11796 7744
rect 10652 7704 11796 7732
rect 10652 7692 10658 7704
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 13262 7692 13268 7744
rect 13320 7692 13326 7744
rect 1104 7642 14904 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 14904 7642
rect 1104 7568 14904 7590
rect 2746 7500 7788 7528
rect 2041 7463 2099 7469
rect 2041 7429 2053 7463
rect 2087 7460 2099 7463
rect 2746 7460 2774 7500
rect 2087 7432 2774 7460
rect 3513 7463 3571 7469
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 3513 7429 3525 7463
rect 3559 7460 3571 7463
rect 3559 7432 3924 7460
rect 3559 7429 3571 7432
rect 3513 7423 3571 7429
rect 3896 7404 3924 7432
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 4028 7432 4077 7460
rect 4028 7420 4034 7432
rect 4065 7429 4077 7432
rect 4111 7460 4123 7463
rect 5258 7460 5264 7472
rect 4111 7432 5264 7460
rect 4111 7429 4123 7432
rect 4065 7423 4123 7429
rect 5258 7420 5264 7432
rect 5316 7460 5322 7472
rect 5442 7460 5448 7472
rect 5316 7432 5448 7460
rect 5316 7420 5322 7432
rect 5442 7420 5448 7432
rect 5500 7460 5506 7472
rect 6454 7460 6460 7472
rect 5500 7432 6460 7460
rect 5500 7420 5506 7432
rect 6454 7420 6460 7432
rect 6512 7420 6518 7472
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3418 7392 3424 7404
rect 3099 7364 3424 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3620 7268 3648 7355
rect 3694 7352 3700 7404
rect 3752 7352 3758 7404
rect 3878 7352 3884 7404
rect 3936 7352 3942 7404
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4614 7392 4620 7404
rect 4295 7364 4620 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 3712 7324 3740 7352
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 3712 7296 3985 7324
rect 3973 7293 3985 7296
rect 4019 7293 4031 7327
rect 6564 7324 6592 7352
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6564 7296 6653 7324
rect 3973 7287 4031 7293
rect 6641 7293 6653 7296
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 3602 7216 3608 7268
rect 3660 7256 3666 7268
rect 4706 7256 4712 7268
rect 3660 7228 4712 7256
rect 3660 7216 3666 7228
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 6748 7256 6776 7355
rect 7760 7324 7788 7500
rect 7834 7488 7840 7540
rect 7892 7488 7898 7540
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 8573 7531 8631 7537
rect 8573 7497 8585 7531
rect 8619 7497 8631 7531
rect 8573 7491 8631 7497
rect 7852 7392 7880 7488
rect 7944 7460 7972 7488
rect 8113 7463 8171 7469
rect 8113 7460 8125 7463
rect 7944 7432 8125 7460
rect 8113 7429 8125 7432
rect 8159 7429 8171 7463
rect 8588 7460 8616 7491
rect 8754 7488 8760 7540
rect 8812 7488 8818 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9493 7531 9551 7537
rect 9493 7528 9505 7531
rect 9180 7500 9505 7528
rect 9180 7488 9186 7500
rect 9493 7497 9505 7500
rect 9539 7497 9551 7531
rect 9493 7491 9551 7497
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10192 7500 11928 7528
rect 10192 7488 10198 7500
rect 9398 7460 9404 7472
rect 8588 7432 9404 7460
rect 8113 7423 8171 7429
rect 9398 7420 9404 7432
rect 9456 7420 9462 7472
rect 11238 7460 11244 7472
rect 9784 7432 11244 7460
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 7852 7364 8677 7392
rect 8665 7361 8677 7364
rect 8711 7392 8723 7395
rect 8846 7392 8852 7404
rect 8711 7364 8852 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9030 7392 9036 7404
rect 8987 7364 9036 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9784 7324 9812 7432
rect 11238 7420 11244 7432
rect 11296 7460 11302 7472
rect 11422 7460 11428 7472
rect 11296 7432 11428 7460
rect 11296 7420 11302 7432
rect 11422 7420 11428 7432
rect 11480 7460 11486 7472
rect 11900 7469 11928 7500
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 11480 7432 11805 7460
rect 11480 7420 11486 7432
rect 11793 7429 11805 7432
rect 11839 7429 11851 7463
rect 11793 7423 11851 7429
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7429 11943 7463
rect 11885 7423 11943 7429
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10410 7392 10416 7404
rect 9907 7364 10416 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10410 7352 10416 7364
rect 10468 7392 10474 7404
rect 10778 7392 10784 7404
rect 10468 7364 10784 7392
rect 10468 7352 10474 7364
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 10870 7352 10876 7404
rect 10928 7352 10934 7404
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11204 7364 11713 7392
rect 11204 7352 11210 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 12032 7364 12081 7392
rect 12032 7352 12038 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 7760 7296 9812 7324
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7324 10011 7327
rect 10226 7324 10232 7336
rect 9999 7296 10232 7324
rect 9999 7293 10011 7296
rect 9953 7287 10011 7293
rect 10226 7284 10232 7296
rect 10284 7324 10290 7336
rect 10888 7324 10916 7352
rect 10284 7296 10916 7324
rect 10284 7284 10290 7296
rect 11514 7284 11520 7336
rect 11572 7284 11578 7336
rect 6656 7228 6776 7256
rect 8481 7259 8539 7265
rect 6656 7200 6684 7228
rect 8481 7225 8493 7259
rect 8527 7256 8539 7259
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 8527 7228 9137 7256
rect 8527 7225 8539 7228
rect 8481 7219 8539 7225
rect 9125 7225 9137 7228
rect 9171 7256 9183 7259
rect 9171 7228 10732 7256
rect 9171 7225 9183 7228
rect 9125 7219 9183 7225
rect 10704 7200 10732 7228
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 5258 7188 5264 7200
rect 4488 7160 5264 7188
rect 4488 7148 4494 7160
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 6638 7148 6644 7200
rect 6696 7148 6702 7200
rect 6733 7191 6791 7197
rect 6733 7157 6745 7191
rect 6779 7188 6791 7191
rect 6822 7188 6828 7200
rect 6779 7160 6828 7188
rect 6779 7157 6791 7160
rect 6733 7151 6791 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 6917 7191 6975 7197
rect 6917 7157 6929 7191
rect 6963 7188 6975 7191
rect 7006 7188 7012 7200
rect 6963 7160 7012 7188
rect 6963 7157 6975 7160
rect 6917 7151 6975 7157
rect 7006 7148 7012 7160
rect 7064 7188 7070 7200
rect 8386 7188 8392 7200
rect 7064 7160 8392 7188
rect 7064 7148 7070 7160
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10137 7191 10195 7197
rect 10137 7188 10149 7191
rect 9732 7160 10149 7188
rect 9732 7148 9738 7160
rect 10137 7157 10149 7160
rect 10183 7157 10195 7191
rect 10137 7151 10195 7157
rect 10686 7148 10692 7200
rect 10744 7148 10750 7200
rect 11532 7197 11560 7284
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 1104 7098 14904 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 14214 7098
rect 14266 7046 14278 7098
rect 14330 7046 14342 7098
rect 14394 7046 14406 7098
rect 14458 7046 14470 7098
rect 14522 7046 14904 7098
rect 1104 7024 14904 7046
rect 4157 6987 4215 6993
rect 4157 6984 4169 6987
rect 3344 6956 4169 6984
rect 2866 6740 2872 6792
rect 2924 6780 2930 6792
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2924 6752 2973 6780
rect 2924 6740 2930 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3142 6740 3148 6792
rect 3200 6740 3206 6792
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3344 6789 3372 6956
rect 4157 6953 4169 6956
rect 4203 6953 4215 6987
rect 4157 6947 4215 6953
rect 4341 6987 4399 6993
rect 4341 6953 4353 6987
rect 4387 6984 4399 6987
rect 4614 6984 4620 6996
rect 4387 6956 4620 6984
rect 4387 6953 4399 6956
rect 4341 6947 4399 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 4985 6987 5043 6993
rect 4985 6953 4997 6987
rect 5031 6953 5043 6987
rect 4985 6947 5043 6953
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 5718 6984 5724 6996
rect 5215 6956 5724 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 3513 6919 3571 6925
rect 3513 6885 3525 6919
rect 3559 6916 3571 6919
rect 3602 6916 3608 6928
rect 3559 6888 3608 6916
rect 3559 6885 3571 6888
rect 3513 6879 3571 6885
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 4798 6916 4804 6928
rect 4172 6888 4804 6916
rect 3786 6808 3792 6860
rect 3844 6808 3850 6860
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 3292 6752 3341 6780
rect 3292 6740 3298 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 4062 6780 4068 6792
rect 3568 6752 4068 6780
rect 3568 6740 3574 6752
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 4172 6721 4200 6888
rect 4798 6876 4804 6888
rect 4856 6916 4862 6928
rect 5000 6916 5028 6947
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 5813 6987 5871 6993
rect 5813 6953 5825 6987
rect 5859 6984 5871 6987
rect 5859 6956 6224 6984
rect 5859 6953 5871 6956
rect 5813 6947 5871 6953
rect 4856 6888 5028 6916
rect 4856 6876 4862 6888
rect 4246 6808 4252 6860
rect 4304 6808 4310 6860
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 4706 6848 4712 6860
rect 4663 6820 4712 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 4706 6808 4712 6820
rect 4764 6848 4770 6860
rect 5828 6848 5856 6947
rect 6196 6925 6224 6956
rect 8938 6944 8944 6996
rect 8996 6984 9002 6996
rect 10870 6984 10876 6996
rect 8996 6956 10876 6984
rect 8996 6944 9002 6956
rect 10870 6944 10876 6956
rect 10928 6984 10934 6996
rect 11698 6984 11704 6996
rect 10928 6956 11704 6984
rect 10928 6944 10934 6956
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 6181 6919 6239 6925
rect 6181 6885 6193 6919
rect 6227 6916 6239 6919
rect 6822 6916 6828 6928
rect 6227 6888 6828 6916
rect 6227 6885 6239 6888
rect 6181 6879 6239 6885
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 10597 6919 10655 6925
rect 10597 6885 10609 6919
rect 10643 6885 10655 6919
rect 10597 6879 10655 6885
rect 4764 6820 5856 6848
rect 4764 6808 4770 6820
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 8570 6848 8576 6860
rect 5960 6820 8576 6848
rect 5960 6808 5966 6820
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 8987 6820 9597 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6848 9827 6851
rect 10612 6848 10640 6879
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 10744 6888 11836 6916
rect 10744 6876 10750 6888
rect 11808 6848 11836 6888
rect 12713 6851 12771 6857
rect 9815 6820 10548 6848
rect 10612 6820 11744 6848
rect 11808 6820 12434 6848
rect 9815 6817 9827 6820
rect 9769 6811 9827 6817
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 3099 6684 4169 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 4157 6681 4169 6684
rect 4203 6681 4215 6715
rect 4264 6712 4292 6808
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 4890 6780 4896 6792
rect 4580 6752 4896 6780
rect 4580 6740 4586 6752
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 5000 6752 5672 6780
rect 5000 6721 5028 6752
rect 4985 6715 5043 6721
rect 4985 6712 4997 6715
rect 4264 6684 4997 6712
rect 4157 6675 4215 6681
rect 4985 6681 4997 6684
rect 5031 6681 5043 6715
rect 4985 6675 5043 6681
rect 5353 6715 5411 6721
rect 5353 6681 5365 6715
rect 5399 6712 5411 6715
rect 5442 6712 5448 6724
rect 5399 6684 5448 6712
rect 5399 6681 5411 6684
rect 5353 6675 5411 6681
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 5644 6712 5672 6752
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6638 6780 6644 6792
rect 5859 6752 6644 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 5828 6712 5856 6743
rect 6638 6740 6644 6752
rect 6696 6780 6702 6792
rect 6733 6783 6791 6789
rect 6733 6780 6745 6783
rect 6696 6752 6745 6780
rect 6696 6740 6702 6752
rect 6733 6749 6745 6752
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8536 6752 9137 6780
rect 8536 6740 8542 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 5644 6684 5856 6712
rect 5920 6684 6193 6712
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 5920 6644 5948 6684
rect 6181 6681 6193 6684
rect 6227 6712 6239 6715
rect 6454 6712 6460 6724
rect 6227 6684 6460 6712
rect 6227 6681 6239 6684
rect 6181 6675 6239 6681
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 5776 6616 5948 6644
rect 5776 6604 5782 6616
rect 5994 6604 6000 6656
rect 6052 6604 6058 6656
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 6420 6616 6653 6644
rect 6420 6604 6426 6616
rect 6641 6613 6653 6616
rect 6687 6613 6699 6647
rect 6641 6607 6699 6613
rect 6914 6604 6920 6656
rect 6972 6604 6978 6656
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 9272 6616 9321 6644
rect 9272 6604 9278 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 9416 6644 9444 6743
rect 9508 6712 9536 6743
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9732 6752 9873 6780
rect 9732 6740 9738 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 9953 6715 10011 6721
rect 9953 6712 9965 6715
rect 9508 6684 9965 6712
rect 9953 6681 9965 6684
rect 9999 6681 10011 6715
rect 9953 6675 10011 6681
rect 9674 6644 9680 6656
rect 9416 6616 9680 6644
rect 9309 6607 9367 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9766 6604 9772 6656
rect 9824 6604 9830 6656
rect 9858 6604 9864 6656
rect 9916 6644 9922 6656
rect 10060 6644 10088 6743
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 10192 6752 10333 6780
rect 10192 6740 10198 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10336 6712 10364 6743
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10336 6684 10456 6712
rect 10428 6656 10456 6684
rect 9916 6616 10088 6644
rect 9916 6604 9922 6616
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 10520 6644 10548 6820
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 10870 6740 10876 6792
rect 10928 6740 10934 6792
rect 10962 6740 10968 6792
rect 11020 6740 11026 6792
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 11103 6752 11192 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 10594 6672 10600 6724
rect 10652 6672 10658 6724
rect 11164 6712 11192 6752
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6780 11483 6783
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11471 6752 11529 6780
rect 11471 6749 11483 6752
rect 11425 6743 11483 6749
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11606 6740 11612 6792
rect 11664 6740 11670 6792
rect 11716 6789 11744 6820
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11624 6712 11652 6740
rect 11164 6684 11652 6712
rect 11808 6712 11836 6743
rect 11882 6740 11888 6792
rect 11940 6740 11946 6792
rect 12406 6712 12434 6820
rect 12713 6817 12725 6851
rect 12759 6848 12771 6851
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12759 6820 12909 6848
rect 12759 6817 12771 6820
rect 12713 6811 12771 6817
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13096 6712 13124 6743
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 11808 6684 12296 6712
rect 12406 6684 13124 6712
rect 12268 6653 12296 6684
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 10520 6616 12173 6644
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 12253 6647 12311 6653
rect 12253 6613 12265 6647
rect 12299 6613 12311 6647
rect 12253 6607 12311 6613
rect 1104 6554 14904 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 14904 6554
rect 1104 6480 14904 6502
rect 3789 6443 3847 6449
rect 3789 6409 3801 6443
rect 3835 6440 3847 6443
rect 3878 6440 3884 6452
rect 3835 6412 3884 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 2777 6375 2835 6381
rect 2777 6341 2789 6375
rect 2823 6372 2835 6375
rect 3804 6372 3832 6403
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 4304 6412 4660 6440
rect 4304 6400 4310 6412
rect 2823 6344 3832 6372
rect 2823 6341 2835 6344
rect 2777 6335 2835 6341
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 4522 6332 4528 6384
rect 4580 6332 4586 6384
rect 4632 6381 4660 6412
rect 4798 6400 4804 6452
rect 4856 6400 4862 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5534 6440 5540 6452
rect 5031 6412 5540 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 7006 6440 7012 6452
rect 6696 6412 7012 6440
rect 6696 6400 6702 6412
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7561 6443 7619 6449
rect 7561 6440 7573 6443
rect 7156 6412 7573 6440
rect 7156 6400 7162 6412
rect 7561 6409 7573 6412
rect 7607 6409 7619 6443
rect 7561 6403 7619 6409
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10686 6440 10692 6452
rect 10643 6412 10692 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 10962 6400 10968 6452
rect 11020 6440 11026 6452
rect 11146 6440 11152 6452
rect 11020 6412 11152 6440
rect 11020 6400 11026 6412
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 12618 6440 12624 6452
rect 12406 6412 12624 6440
rect 4617 6375 4675 6381
rect 4617 6341 4629 6375
rect 4663 6341 4675 6375
rect 6012 6372 6040 6400
rect 9858 6372 9864 6384
rect 6012 6344 7144 6372
rect 4617 6335 4675 6341
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3418 6304 3424 6316
rect 3283 6276 3424 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6304 3571 6307
rect 3988 6304 4016 6332
rect 3559 6276 4016 6304
rect 4249 6307 4307 6313
rect 3559 6273 3571 6276
rect 3513 6267 3571 6273
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4540 6304 4568 6332
rect 4295 6276 4568 6304
rect 6549 6307 6607 6313
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 6914 6304 6920 6316
rect 6687 6276 6920 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3326 6236 3332 6248
rect 3191 6208 3332 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3326 6196 3332 6208
rect 3384 6236 3390 6248
rect 3528 6236 3556 6267
rect 3384 6208 3556 6236
rect 3881 6239 3939 6245
rect 3384 6196 3390 6208
rect 3881 6205 3893 6239
rect 3927 6205 3939 6239
rect 3881 6199 3939 6205
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 3896 6168 3924 6199
rect 3252 6140 3924 6168
rect 3252 6112 3280 6140
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 3234 6100 3240 6112
rect 2924 6072 3240 6100
rect 2924 6060 2930 6072
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 3418 6060 3424 6112
rect 3476 6060 3482 6112
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 3988 6100 4016 6199
rect 6564 6180 6592 6267
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 7116 6313 7144 6344
rect 8772 6344 8984 6372
rect 8772 6316 8800 6344
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8754 6304 8760 6316
rect 8619 6276 8760 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6205 7895 6239
rect 7837 6199 7895 6205
rect 6546 6128 6552 6180
rect 6604 6168 6610 6180
rect 7852 6168 7880 6199
rect 7926 6196 7932 6248
rect 7984 6236 7990 6248
rect 8128 6236 8156 6267
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 8956 6313 8984 6344
rect 9232 6344 9864 6372
rect 9232 6316 9260 6344
rect 9858 6332 9864 6344
rect 9916 6372 9922 6384
rect 12406 6372 12434 6412
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 12897 6443 12955 6449
rect 12897 6409 12909 6443
rect 12943 6440 12955 6443
rect 13354 6440 13360 6452
rect 12943 6412 13360 6440
rect 12943 6409 12955 6412
rect 12897 6403 12955 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 9916 6344 12434 6372
rect 9916 6332 9922 6344
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 9088 6276 9137 6304
rect 9088 6264 9094 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9214 6264 9220 6316
rect 9272 6264 9278 6316
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10502 6304 10508 6316
rect 10459 6276 10508 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 7984 6208 8800 6236
rect 7984 6196 7990 6208
rect 6604 6140 7880 6168
rect 6604 6128 6610 6140
rect 3844 6072 4016 6100
rect 3844 6060 3850 6072
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4764 6072 4813 6100
rect 4764 6060 4770 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8665 6103 8723 6109
rect 8665 6100 8677 6103
rect 8260 6072 8677 6100
rect 8260 6060 8266 6072
rect 8665 6069 8677 6072
rect 8711 6069 8723 6103
rect 8772 6100 8800 6208
rect 8846 6128 8852 6180
rect 8904 6168 8910 6180
rect 9324 6168 9352 6267
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10778 6304 10784 6316
rect 10643 6276 10784 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 11900 6236 11928 6264
rect 9456 6208 11928 6236
rect 9456 6196 9462 6208
rect 12406 6180 12434 6344
rect 12802 6264 12808 6316
rect 12860 6264 12866 6316
rect 14461 6307 14519 6313
rect 14461 6273 14473 6307
rect 14507 6304 14519 6307
rect 14918 6304 14924 6316
rect 14507 6276 14924 6304
rect 14507 6273 14519 6276
rect 14461 6267 14519 6273
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 8904 6140 9352 6168
rect 9769 6171 9827 6177
rect 8904 6128 8910 6140
rect 9769 6137 9781 6171
rect 9815 6137 9827 6171
rect 12406 6140 12440 6180
rect 9769 6131 9827 6137
rect 9401 6103 9459 6109
rect 9401 6100 9413 6103
rect 8772 6072 9413 6100
rect 8665 6063 8723 6069
rect 9401 6069 9413 6072
rect 9447 6069 9459 6103
rect 9401 6063 9459 6069
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 9784 6100 9812 6131
rect 12434 6128 12440 6140
rect 12492 6128 12498 6180
rect 9640 6072 9812 6100
rect 9640 6060 9646 6072
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 11112 6072 14381 6100
rect 11112 6060 11118 6072
rect 14369 6069 14381 6072
rect 14415 6069 14427 6103
rect 14369 6063 14427 6069
rect 1104 6010 14904 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 14214 6010
rect 14266 5958 14278 6010
rect 14330 5958 14342 6010
rect 14394 5958 14406 6010
rect 14458 5958 14470 6010
rect 14522 5958 14904 6010
rect 1104 5936 14904 5958
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3384 5868 3433 5896
rect 3384 5856 3390 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 3421 5859 3479 5865
rect 5350 5856 5356 5908
rect 5408 5856 5414 5908
rect 7006 5856 7012 5908
rect 7064 5856 7070 5908
rect 7926 5856 7932 5908
rect 7984 5856 7990 5908
rect 8113 5899 8171 5905
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 9030 5896 9036 5908
rect 8159 5868 9036 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9582 5856 9588 5908
rect 9640 5856 9646 5908
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 11149 5899 11207 5905
rect 11149 5896 11161 5899
rect 10652 5868 11161 5896
rect 10652 5856 10658 5868
rect 11149 5865 11161 5868
rect 11195 5865 11207 5899
rect 11149 5859 11207 5865
rect 12434 5856 12440 5908
rect 12492 5856 12498 5908
rect 9600 5828 9628 5856
rect 7944 5800 9628 5828
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 4798 5760 4804 5772
rect 2188 5732 4804 5760
rect 2188 5720 2194 5732
rect 4798 5720 4804 5732
rect 4856 5760 4862 5772
rect 5537 5763 5595 5769
rect 4856 5732 5120 5760
rect 4856 5720 4862 5732
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 5092 5701 5120 5732
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 5583 5732 6837 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3476 5664 3801 5692
rect 3476 5652 3482 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 7834 5692 7840 5704
rect 6779 5664 7840 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 3142 5584 3148 5636
rect 3200 5624 3206 5636
rect 3513 5627 3571 5633
rect 3513 5624 3525 5627
rect 3200 5596 3525 5624
rect 3200 5584 3206 5596
rect 3513 5593 3525 5596
rect 3559 5624 3571 5627
rect 6656 5624 6684 5655
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 7944 5624 7972 5800
rect 10318 5788 10324 5840
rect 10376 5828 10382 5840
rect 12802 5828 12808 5840
rect 10376 5800 12808 5828
rect 10376 5788 10382 5800
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 9214 5760 9220 5772
rect 8067 5732 9220 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 13814 5760 13820 5772
rect 9324 5732 13820 5760
rect 8242 5695 8300 5701
rect 8242 5692 8254 5695
rect 8036 5664 8254 5692
rect 8036 5636 8064 5664
rect 8242 5661 8254 5664
rect 8288 5661 8300 5695
rect 8242 5655 8300 5661
rect 3559 5596 6408 5624
rect 6656 5596 7972 5624
rect 3559 5593 3571 5596
rect 3513 5587 3571 5593
rect 3970 5516 3976 5568
rect 4028 5516 4034 5568
rect 6380 5556 6408 5596
rect 8018 5584 8024 5636
rect 8076 5584 8082 5636
rect 8386 5584 8392 5636
rect 8444 5584 8450 5636
rect 9324 5556 9352 5732
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 11330 5701 11336 5704
rect 11309 5695 11336 5701
rect 11309 5661 11321 5695
rect 11309 5655 11336 5661
rect 11330 5652 11336 5655
rect 11388 5652 11394 5704
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 11790 5692 11796 5704
rect 11747 5664 11796 5692
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 12526 5652 12532 5704
rect 12584 5652 12590 5704
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 11425 5627 11483 5633
rect 11425 5624 11437 5627
rect 10652 5596 11437 5624
rect 10652 5584 10658 5596
rect 11425 5593 11437 5596
rect 11471 5593 11483 5627
rect 11425 5587 11483 5593
rect 11514 5584 11520 5636
rect 11572 5584 11578 5636
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 12492 5596 12725 5624
rect 12492 5584 12498 5596
rect 12713 5593 12725 5596
rect 12759 5593 12771 5627
rect 12713 5587 12771 5593
rect 6380 5528 9352 5556
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 11054 5556 11060 5568
rect 9456 5528 11060 5556
rect 9456 5516 9462 5528
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 1104 5466 14904 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 14904 5466
rect 1104 5392 14904 5414
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 5810 5352 5816 5364
rect 5583 5324 5816 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 5810 5312 5816 5324
rect 5868 5352 5874 5364
rect 6822 5352 6828 5364
rect 5868 5324 6500 5352
rect 5868 5312 5874 5324
rect 4724 5256 5304 5284
rect 4724 5225 4752 5256
rect 5276 5228 5304 5256
rect 5350 5244 5356 5296
rect 5408 5284 5414 5296
rect 6472 5293 6500 5324
rect 6748 5324 6828 5352
rect 6457 5287 6515 5293
rect 5408 5256 5856 5284
rect 5408 5244 5414 5256
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4856 5188 5181 5216
rect 4856 5176 4862 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5258 5176 5264 5228
rect 5316 5176 5322 5228
rect 5442 5176 5448 5228
rect 5500 5216 5506 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5500 5188 5641 5216
rect 5500 5176 5506 5188
rect 5629 5185 5641 5188
rect 5675 5216 5687 5219
rect 5718 5216 5724 5228
rect 5675 5188 5724 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 5828 5225 5856 5256
rect 6457 5253 6469 5287
rect 6503 5253 6515 5287
rect 6457 5247 6515 5253
rect 6748 5225 6776 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 8113 5355 8171 5361
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 8159 5324 8432 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8404 5296 8432 5324
rect 9508 5324 11008 5352
rect 8202 5284 8208 5296
rect 7944 5256 8208 5284
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 6733 5219 6791 5225
rect 5859 5188 6500 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 4893 5151 4951 5157
rect 4893 5117 4905 5151
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5031 5120 5488 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 4908 5080 4936 5111
rect 5350 5080 5356 5092
rect 4908 5052 5356 5080
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 4614 5012 4620 5024
rect 4571 4984 4620 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 5460 5012 5488 5120
rect 6362 5108 6368 5160
rect 6420 5108 6426 5160
rect 6472 5148 6500 5188
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7006 5216 7012 5228
rect 6871 5188 7012 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7944 5225 7972 5256
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 8386 5244 8392 5296
rect 8444 5244 8450 5296
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5185 7987 5219
rect 7929 5179 7987 5185
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 8110 5216 8116 5228
rect 8067 5188 8116 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 8110 5176 8116 5188
rect 8168 5216 8174 5228
rect 9508 5216 9536 5324
rect 10152 5256 10732 5284
rect 8168 5188 9536 5216
rect 9585 5219 9643 5225
rect 8168 5176 8174 5188
rect 9585 5185 9597 5219
rect 9631 5216 9643 5219
rect 9950 5216 9956 5228
rect 9631 5188 9956 5216
rect 9631 5185 9643 5188
rect 9585 5179 9643 5185
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10152 5225 10180 5256
rect 10704 5228 10732 5256
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10284 5188 10425 5216
rect 10284 5176 10290 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 10502 5176 10508 5228
rect 10560 5176 10566 5228
rect 10594 5176 10600 5228
rect 10652 5176 10658 5228
rect 10686 5176 10692 5228
rect 10744 5176 10750 5228
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 8297 5151 8355 5157
rect 6472 5120 8230 5148
rect 8202 5080 8230 5120
rect 8297 5117 8309 5151
rect 8343 5148 8355 5151
rect 8478 5148 8484 5160
rect 8343 5120 8484 5148
rect 8343 5117 8355 5120
rect 8297 5111 8355 5117
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 9398 5108 9404 5160
rect 9456 5108 9462 5160
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5117 9735 5151
rect 9677 5111 9735 5117
rect 9416 5080 9444 5108
rect 8202 5052 9444 5080
rect 9692 5080 9720 5111
rect 10042 5108 10048 5160
rect 10100 5108 10106 5160
rect 10318 5108 10324 5160
rect 10376 5108 10382 5160
rect 10612 5148 10640 5176
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 10612 5120 10793 5148
rect 10781 5117 10793 5120
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 10137 5083 10195 5089
rect 10137 5080 10149 5083
rect 9692 5052 10149 5080
rect 10137 5049 10149 5052
rect 10183 5049 10195 5083
rect 10888 5080 10916 5179
rect 10137 5043 10195 5049
rect 10244 5052 10916 5080
rect 10980 5080 11008 5324
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 12345 5355 12403 5361
rect 12345 5352 12357 5355
rect 11204 5324 12357 5352
rect 11204 5312 11210 5324
rect 12345 5321 12357 5324
rect 12391 5321 12403 5355
rect 12345 5315 12403 5321
rect 12434 5312 12440 5364
rect 12492 5312 12498 5364
rect 13354 5312 13360 5364
rect 13412 5312 13418 5364
rect 11238 5244 11244 5296
rect 11296 5244 11302 5296
rect 12452 5284 12480 5312
rect 13372 5284 13400 5312
rect 12268 5256 12940 5284
rect 12268 5225 12296 5256
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 12526 5216 12532 5228
rect 12483 5188 12532 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 11146 5108 11152 5160
rect 11204 5108 11210 5160
rect 12912 5148 12940 5256
rect 13004 5256 13400 5284
rect 13004 5225 13032 5256
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 13127 5188 13185 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13449 5219 13507 5225
rect 13449 5185 13461 5219
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 13096 5148 13124 5179
rect 12912 5120 13124 5148
rect 13262 5080 13268 5092
rect 10980 5052 12434 5080
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 5460 4984 5641 5012
rect 5629 4981 5641 4984
rect 5675 4981 5687 5015
rect 5629 4975 5687 4981
rect 7006 4972 7012 5024
rect 7064 4972 7070 5024
rect 8018 4972 8024 5024
rect 8076 4972 8082 5024
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 9180 4984 9413 5012
rect 9180 4972 9186 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 9401 4975 9459 4981
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10244 5012 10272 5052
rect 9640 4984 10272 5012
rect 9640 4972 9646 4984
rect 10318 4972 10324 5024
rect 10376 5012 10382 5024
rect 10597 5015 10655 5021
rect 10597 5012 10609 5015
rect 10376 4984 10609 5012
rect 10376 4972 10382 4984
rect 10597 4981 10609 4984
rect 10643 4981 10655 5015
rect 10888 5012 10916 5052
rect 11606 5012 11612 5024
rect 10888 4984 11612 5012
rect 10597 4975 10655 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 12406 5012 12434 5052
rect 13096 5052 13268 5080
rect 13096 5021 13124 5052
rect 13262 5040 13268 5052
rect 13320 5080 13326 5092
rect 13464 5080 13492 5179
rect 13320 5052 13492 5080
rect 13320 5040 13326 5052
rect 12713 5015 12771 5021
rect 12713 5012 12725 5015
rect 12406 4984 12725 5012
rect 12713 4981 12725 4984
rect 12759 4981 12771 5015
rect 12713 4975 12771 4981
rect 13081 5015 13139 5021
rect 13081 4981 13093 5015
rect 13127 4981 13139 5015
rect 13081 4975 13139 4981
rect 13170 4972 13176 5024
rect 13228 4972 13234 5024
rect 1104 4922 14904 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 14214 4922
rect 14266 4870 14278 4922
rect 14330 4870 14342 4922
rect 14394 4870 14406 4922
rect 14458 4870 14470 4922
rect 14522 4870 14904 4922
rect 1104 4848 14904 4870
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 6641 4811 6699 4817
rect 6641 4808 6653 4811
rect 6420 4780 6653 4808
rect 6420 4768 6426 4780
rect 6641 4777 6653 4780
rect 6687 4777 6699 4811
rect 6641 4771 6699 4777
rect 7101 4811 7159 4817
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 7650 4808 7656 4820
rect 7147 4780 7656 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 7650 4768 7656 4780
rect 7708 4808 7714 4820
rect 7926 4808 7932 4820
rect 7708 4780 7932 4808
rect 7708 4768 7714 4780
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8018 4768 8024 4820
rect 8076 4768 8082 4820
rect 11241 4811 11299 4817
rect 11241 4777 11253 4811
rect 11287 4808 11299 4811
rect 11514 4808 11520 4820
rect 11287 4780 11520 4808
rect 11287 4777 11299 4780
rect 11241 4771 11299 4777
rect 5810 4700 5816 4752
rect 5868 4740 5874 4752
rect 6822 4740 6828 4752
rect 5868 4712 6828 4740
rect 5868 4700 5874 4712
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 7742 4700 7748 4752
rect 7800 4740 7806 4752
rect 7837 4743 7895 4749
rect 7837 4740 7849 4743
rect 7800 4712 7849 4740
rect 7800 4700 7806 4712
rect 7837 4709 7849 4712
rect 7883 4709 7895 4743
rect 8036 4740 8064 4768
rect 10686 4740 10692 4752
rect 8036 4712 8156 4740
rect 7837 4703 7895 4709
rect 8128 4681 8156 4712
rect 9784 4712 10692 4740
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 5552 4644 6469 4672
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4856 4576 4997 4604
rect 4856 4564 4862 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5350 4604 5356 4616
rect 5215 4576 5356 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5552 4480 5580 4644
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 6380 4594 6408 4644
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 8113 4675 8171 4681
rect 8113 4641 8125 4675
rect 8159 4641 8171 4675
rect 8113 4635 8171 4641
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 8570 4672 8576 4684
rect 8251 4644 8576 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 6288 4536 6316 4567
rect 6380 4566 6592 4594
rect 6564 4536 6592 4566
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4606 6791 4607
rect 6822 4606 6828 4616
rect 6779 4578 6828 4606
rect 6779 4573 6791 4578
rect 6733 4567 6791 4573
rect 6822 4564 6828 4578
rect 6880 4564 6886 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 6932 4536 6960 4567
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7800 4576 8033 4604
rect 7800 4564 7806 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 6288 4508 6500 4536
rect 6564 4508 6960 4536
rect 9600 4536 9628 4567
rect 9674 4564 9680 4616
rect 9732 4564 9738 4616
rect 9784 4604 9812 4712
rect 10686 4700 10692 4712
rect 10744 4740 10750 4752
rect 11256 4740 11284 4771
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 12434 4808 12440 4820
rect 12299 4780 12440 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 13872 4780 14381 4808
rect 13872 4768 13878 4780
rect 14369 4777 14381 4780
rect 14415 4777 14427 4811
rect 14369 4771 14427 4777
rect 10744 4712 11284 4740
rect 10744 4700 10750 4712
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 12345 4743 12403 4749
rect 12345 4740 12357 4743
rect 11480 4712 12357 4740
rect 11480 4700 11486 4712
rect 12345 4709 12357 4712
rect 12391 4709 12403 4743
rect 12345 4703 12403 4709
rect 11440 4644 11744 4672
rect 9846 4607 9904 4613
rect 9846 4604 9858 4607
rect 9784 4576 9858 4604
rect 9846 4573 9858 4576
rect 9892 4573 9904 4607
rect 9846 4567 9904 4573
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 10042 4604 10048 4616
rect 9999 4576 10048 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 11440 4613 11468 4644
rect 11716 4616 11744 4644
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 11514 4564 11520 4616
rect 11572 4564 11578 4616
rect 11698 4564 11704 4616
rect 11756 4604 11762 4616
rect 12069 4607 12127 4613
rect 12069 4604 12081 4607
rect 11756 4576 12081 4604
rect 11756 4564 11762 4576
rect 12069 4573 12081 4576
rect 12115 4604 12127 4607
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12115 4576 12725 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4604 14611 4607
rect 14599 4576 14964 4604
rect 14599 4573 14611 4576
rect 14553 4567 14611 4573
rect 11532 4536 11560 4564
rect 11885 4539 11943 4545
rect 11885 4536 11897 4539
rect 9600 4508 10548 4536
rect 11532 4508 11897 4536
rect 6472 4480 6500 4508
rect 10520 4480 10548 4508
rect 11885 4505 11897 4508
rect 11931 4505 11943 4539
rect 11885 4499 11943 4505
rect 14936 4480 14964 4576
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 4798 4468 4804 4480
rect 1627 4440 4804 4468
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4468 5227 4471
rect 5534 4468 5540 4480
rect 5215 4440 5540 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 6362 4428 6368 4480
rect 6420 4428 6426 4480
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 6914 4468 6920 4480
rect 6512 4440 6920 4468
rect 6512 4428 6518 4440
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 9030 4468 9036 4480
rect 7064 4440 9036 4468
rect 7064 4428 7070 4440
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 9214 4428 9220 4480
rect 9272 4468 9278 4480
rect 9401 4471 9459 4477
rect 9401 4468 9413 4471
rect 9272 4440 9413 4468
rect 9272 4428 9278 4440
rect 9401 4437 9413 4440
rect 9447 4437 9459 4471
rect 9401 4431 9459 4437
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 11701 4471 11759 4477
rect 11701 4468 11713 4471
rect 10560 4440 11713 4468
rect 10560 4428 10566 4440
rect 11701 4437 11713 4440
rect 11747 4437 11759 4471
rect 11701 4431 11759 4437
rect 14918 4428 14924 4480
rect 14976 4428 14982 4480
rect 1104 4378 14904 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 14904 4378
rect 1104 4304 14904 4326
rect 5534 4224 5540 4276
rect 5592 4224 5598 4276
rect 8202 4224 8208 4276
rect 8260 4224 8266 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8352 4236 8953 4264
rect 8352 4224 8358 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 8941 4227 8999 4233
rect 9030 4224 9036 4276
rect 9088 4264 9094 4276
rect 13906 4264 13912 4276
rect 9088 4236 13912 4264
rect 9088 4224 9094 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 5077 4199 5135 4205
rect 5077 4165 5089 4199
rect 5123 4196 5135 4199
rect 5123 4168 5488 4196
rect 5123 4165 5135 4168
rect 5077 4159 5135 4165
rect 4614 4088 4620 4140
rect 4672 4128 4678 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 4672 4100 4721 4128
rect 4672 4088 4678 4100
rect 4709 4097 4721 4100
rect 4755 4097 4767 4131
rect 4709 4091 4767 4097
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 4856 4100 4936 4128
rect 4856 4088 4862 4100
rect 4908 3992 4936 4100
rect 4982 4088 4988 4140
rect 5040 4088 5046 4140
rect 5215 4131 5273 4137
rect 5215 4097 5227 4131
rect 5261 4128 5273 4131
rect 5350 4128 5356 4140
rect 5261 4100 5356 4128
rect 5261 4097 5273 4100
rect 5215 4091 5273 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5460 4137 5488 4168
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4097 5503 4131
rect 5552 4128 5580 4224
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5552 4100 5641 4128
rect 5445 4091 5503 4097
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8220 4128 8248 4224
rect 10318 4196 10324 4208
rect 8159 4100 8248 4128
rect 8680 4168 10088 4196
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 5460 4060 5488 4091
rect 5810 4060 5816 4072
rect 5460 4032 5816 4060
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4029 8355 4063
rect 8297 4023 8355 4029
rect 4908 3964 8064 3992
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 5442 3924 5448 3936
rect 5399 3896 5448 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 7800 3896 7941 3924
rect 7800 3884 7806 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 8036 3924 8064 3964
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 8220 3992 8248 4023
rect 8168 3964 8248 3992
rect 8312 3992 8340 4023
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8680 4060 8708 4168
rect 10060 4140 10088 4168
rect 10244 4168 10324 4196
rect 9122 4088 9128 4140
rect 9180 4088 9186 4140
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 9490 4128 9496 4140
rect 9355 4100 9496 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 9858 4088 9864 4140
rect 9916 4088 9922 4140
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10042 4088 10048 4140
rect 10100 4088 10106 4140
rect 10134 4088 10140 4140
rect 10192 4088 10198 4140
rect 10244 4137 10272 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 11572 4168 12020 4196
rect 11572 4156 11578 4168
rect 11992 4137 12020 4168
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12066 4128 12072 4140
rect 12023 4100 12072 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 8444 4032 8708 4060
rect 8444 4020 8450 4032
rect 9214 4020 9220 4072
rect 9272 4020 9278 4072
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9447 4032 9689 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 8478 3992 8484 4004
rect 8312 3964 8484 3992
rect 8168 3952 8174 3964
rect 8478 3952 8484 3964
rect 8536 3992 8542 4004
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 8536 3964 11529 3992
rect 8536 3952 8542 3964
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 11517 3955 11575 3961
rect 9306 3924 9312 3936
rect 8036 3896 9312 3924
rect 7929 3887 7987 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10778 3924 10784 3936
rect 9732 3896 10784 3924
rect 9732 3884 9738 3896
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 11698 3884 11704 3936
rect 11756 3884 11762 3936
rect 1104 3834 14904 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 14214 3834
rect 14266 3782 14278 3834
rect 14330 3782 14342 3834
rect 14394 3782 14406 3834
rect 14458 3782 14470 3834
rect 14522 3782 14904 3834
rect 1104 3760 14904 3782
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5040 3692 7788 3720
rect 5040 3680 5046 3692
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 6181 3655 6239 3661
rect 6181 3652 6193 3655
rect 5316 3624 6193 3652
rect 5316 3612 5322 3624
rect 6181 3621 6193 3624
rect 6227 3621 6239 3655
rect 6181 3615 6239 3621
rect 6454 3612 6460 3664
rect 6512 3612 6518 3664
rect 6638 3612 6644 3664
rect 6696 3652 6702 3664
rect 6914 3652 6920 3664
rect 6696 3624 6920 3652
rect 6696 3612 6702 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7760 3652 7788 3692
rect 7834 3680 7840 3732
rect 7892 3680 7898 3732
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 8251 3692 9812 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 9784 3652 9812 3692
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9916 3692 9965 3720
rect 9916 3680 9922 3692
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 9953 3683 10011 3689
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10192 3692 10241 3720
rect 10192 3680 10198 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 10229 3683 10287 3689
rect 11790 3680 11796 3732
rect 11848 3680 11854 3732
rect 10318 3652 10324 3664
rect 7760 3624 8294 3652
rect 9784 3624 10324 3652
rect 5902 3544 5908 3596
rect 5960 3544 5966 3596
rect 6086 3476 6092 3528
rect 6144 3476 6150 3528
rect 6362 3476 6368 3528
rect 6420 3476 6426 3528
rect 6472 3525 6500 3612
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7708 3556 8125 3584
rect 7708 3544 7714 3556
rect 8113 3553 8125 3556
rect 8159 3553 8171 3587
rect 8266 3584 8294 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 11808 3652 11836 3680
rect 10428 3624 11836 3652
rect 8266 3556 10272 3584
rect 8113 3547 8171 3553
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 8662 3516 8668 3528
rect 8251 3488 8668 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9732 3488 9781 3516
rect 9732 3476 9738 3488
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 5350 3408 5356 3460
rect 5408 3448 5414 3460
rect 5534 3448 5540 3460
rect 5408 3420 5540 3448
rect 5408 3408 5414 3420
rect 5534 3408 5540 3420
rect 5592 3448 5598 3460
rect 6181 3451 6239 3457
rect 6181 3448 6193 3451
rect 5592 3420 6193 3448
rect 5592 3408 5598 3420
rect 6181 3417 6193 3420
rect 6227 3448 6239 3451
rect 6822 3448 6828 3460
rect 6227 3420 6828 3448
rect 6227 3417 6239 3420
rect 6181 3411 6239 3417
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 9582 3408 9588 3460
rect 9640 3408 9646 3460
rect 4798 3340 4804 3392
rect 4856 3380 4862 3392
rect 8938 3380 8944 3392
rect 4856 3352 8944 3380
rect 4856 3340 4862 3352
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 10244 3380 10272 3556
rect 10428 3525 10456 3624
rect 12066 3612 12072 3664
rect 12124 3612 12130 3664
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 12084 3584 12112 3612
rect 10919 3556 12112 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 10502 3408 10508 3460
rect 10560 3408 10566 3460
rect 10715 3451 10773 3457
rect 10715 3417 10727 3451
rect 10761 3417 10773 3451
rect 10715 3411 10773 3417
rect 10410 3380 10416 3392
rect 10244 3352 10416 3380
rect 10410 3340 10416 3352
rect 10468 3380 10474 3392
rect 10730 3380 10758 3411
rect 11698 3408 11704 3460
rect 11756 3408 11762 3460
rect 10468 3352 10758 3380
rect 12161 3383 12219 3389
rect 10468 3340 10474 3352
rect 12161 3349 12173 3383
rect 12207 3380 12219 3383
rect 12526 3380 12532 3392
rect 12207 3352 12532 3380
rect 12207 3349 12219 3352
rect 12161 3343 12219 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 1104 3290 14904 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 14904 3290
rect 1104 3216 14904 3238
rect 5258 3136 5264 3188
rect 5316 3136 5322 3188
rect 5997 3179 6055 3185
rect 5460 3148 5856 3176
rect 3970 3000 3976 3052
rect 4028 3040 4034 3052
rect 4798 3040 4804 3052
rect 4028 3012 4804 3040
rect 4028 3000 4034 3012
rect 4798 3000 4804 3012
rect 4856 3040 4862 3052
rect 5276 3049 5304 3136
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4856 3012 4997 3040
rect 4856 3000 4862 3012
rect 4985 3009 4997 3012
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5184 2972 5212 3003
rect 5350 3000 5356 3052
rect 5408 3000 5414 3052
rect 5460 3049 5488 3148
rect 5626 3068 5632 3120
rect 5684 3108 5690 3120
rect 5828 3108 5856 3148
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6086 3176 6092 3188
rect 6043 3148 6092 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6457 3179 6515 3185
rect 6457 3145 6469 3179
rect 6503 3145 6515 3179
rect 9401 3179 9459 3185
rect 6457 3139 6515 3145
rect 6748 3148 8892 3176
rect 6472 3108 6500 3139
rect 5684 3080 5764 3108
rect 5828 3080 6500 3108
rect 5684 3068 5690 3080
rect 5736 3049 5764 3080
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 5368 2972 5396 3000
rect 5184 2944 5396 2972
rect 4985 2907 5043 2913
rect 4985 2873 4997 2907
rect 5031 2904 5043 2907
rect 5552 2904 5580 3003
rect 5828 2972 5856 3003
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 6512 3012 6653 3040
rect 6512 3000 6518 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 5031 2876 5580 2904
rect 5736 2944 5856 2972
rect 6380 2972 6408 3000
rect 6748 2981 6776 3148
rect 8570 3108 8576 3120
rect 7300 3080 8432 3108
rect 6914 3000 6920 3052
rect 6972 3000 6978 3052
rect 6733 2975 6791 2981
rect 6733 2972 6745 2975
rect 6380 2944 6745 2972
rect 5031 2873 5043 2876
rect 4985 2867 5043 2873
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5736 2836 5764 2944
rect 6733 2941 6745 2944
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7300 2972 7328 3080
rect 7650 3000 7656 3052
rect 7708 3040 7714 3052
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7708 3012 7757 3040
rect 7708 3000 7714 3012
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 7834 3000 7840 3052
rect 7892 3000 7898 3052
rect 8404 3049 8432 3080
rect 8496 3080 8576 3108
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8389 3043 8447 3049
rect 8159 3012 8340 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 6880 2944 7328 2972
rect 7944 2972 7972 3003
rect 8312 2972 8340 3012
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8496 2972 8524 3080
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 7944 2944 8248 2972
rect 8312 2944 8524 2972
rect 8588 3012 8769 3040
rect 6880 2932 6886 2944
rect 7469 2907 7527 2913
rect 7469 2904 7481 2907
rect 5828 2876 7481 2904
rect 5828 2845 5856 2876
rect 7469 2873 7481 2876
rect 7515 2873 7527 2907
rect 7469 2867 7527 2873
rect 7742 2864 7748 2916
rect 7800 2864 7806 2916
rect 8220 2913 8248 2944
rect 8205 2907 8263 2913
rect 8205 2873 8217 2907
rect 8251 2873 8263 2907
rect 8205 2867 8263 2873
rect 5491 2808 5764 2836
rect 5813 2839 5871 2845
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5813 2805 5825 2839
rect 5859 2805 5871 2839
rect 7760 2836 7788 2864
rect 8588 2836 8616 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8864 2904 8892 3148
rect 9401 3145 9413 3179
rect 9447 3176 9459 3179
rect 9582 3176 9588 3188
rect 9447 3148 9588 3176
rect 9447 3145 9459 3148
rect 9401 3139 9459 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10137 3179 10195 3185
rect 10137 3176 10149 3179
rect 10008 3148 10149 3176
rect 10008 3136 10014 3148
rect 10137 3145 10149 3148
rect 10183 3145 10195 3179
rect 10137 3139 10195 3145
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 10376 3148 12081 3176
rect 10376 3136 10382 3148
rect 12069 3145 12081 3148
rect 12115 3145 12127 3179
rect 12069 3139 12127 3145
rect 8938 3068 8944 3120
rect 8996 3068 9002 3120
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 9968 3040 9996 3136
rect 10042 3068 10048 3120
rect 10100 3068 10106 3120
rect 13170 3108 13176 3120
rect 10336 3080 11560 3108
rect 10336 3049 10364 3080
rect 9907 3012 9996 3040
rect 10321 3043 10379 3049
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10502 3000 10508 3052
rect 10560 3000 10566 3052
rect 10594 3000 10600 3052
rect 10652 3049 10658 3052
rect 10652 3040 10663 3049
rect 10704 3040 10732 3080
rect 10652 3012 10732 3040
rect 10781 3043 10839 3049
rect 10652 3003 10663 3012
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 11054 3040 11060 3052
rect 10827 3012 11060 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 10652 3000 10658 3003
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 9232 2944 9689 2972
rect 9232 2913 9260 2944
rect 9677 2941 9689 2944
rect 9723 2941 9735 2975
rect 10520 2972 10548 3000
rect 10796 2972 10824 3003
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11532 3049 11560 3080
rect 11808 3080 13176 3108
rect 11808 3049 11836 3080
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12526 3040 12532 3052
rect 11931 3012 12532 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 10520 2944 10824 2972
rect 9677 2935 9735 2941
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 8864 2876 9229 2904
rect 9217 2873 9229 2876
rect 9263 2873 9275 2907
rect 9692 2904 9720 2935
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 9692 2876 10701 2904
rect 9217 2867 9275 2873
rect 10689 2873 10701 2876
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 7760 2808 8616 2836
rect 5813 2799 5871 2805
rect 8662 2796 8668 2848
rect 8720 2796 8726 2848
rect 10778 2796 10784 2848
rect 10836 2836 10842 2848
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 10836 2808 10977 2836
rect 10836 2796 10842 2808
rect 10965 2805 10977 2808
rect 11011 2836 11023 2839
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 11011 2808 11621 2836
rect 11011 2805 11023 2808
rect 10965 2799 11023 2805
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 11609 2799 11667 2805
rect 1104 2746 14904 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 14214 2746
rect 14266 2694 14278 2746
rect 14330 2694 14342 2746
rect 14394 2694 14406 2746
rect 14458 2694 14470 2746
rect 14522 2694 14904 2746
rect 1104 2672 14904 2694
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2222 2632 2228 2644
rect 2179 2604 2228 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 2866 2632 2872 2644
rect 2547 2604 2872 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 4157 2635 4215 2641
rect 4157 2632 4169 2635
rect 4120 2604 4169 2632
rect 4120 2592 4126 2604
rect 4157 2601 4169 2604
rect 4203 2601 4215 2635
rect 4157 2595 4215 2601
rect 6178 2592 6184 2644
rect 6236 2592 6242 2644
rect 7653 2635 7711 2641
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 7834 2632 7840 2644
rect 7699 2604 7840 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 11054 2592 11060 2644
rect 11112 2592 11118 2644
rect 1765 2567 1823 2573
rect 1765 2533 1777 2567
rect 1811 2564 1823 2567
rect 6196 2564 6224 2592
rect 1811 2536 6224 2564
rect 1811 2533 1823 2536
rect 1765 2527 1823 2533
rect 7742 2524 7748 2576
rect 7800 2524 7806 2576
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8662 2496 8668 2508
rect 8159 2468 8668 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8662 2456 8668 2468
rect 8720 2496 8726 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8720 2468 8953 2496
rect 8720 2456 8726 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 10778 2496 10784 2508
rect 8941 2459 8999 2465
rect 9140 2468 10784 2496
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 72 2400 1624 2428
rect 72 2388 78 2400
rect 934 2320 940 2372
rect 992 2360 998 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 992 2332 1501 2360
rect 992 2320 998 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1596 2360 1624 2400
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2004 2400 2329 2428
rect 2004 2388 2010 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 6730 2388 6736 2440
rect 6788 2388 6794 2440
rect 9140 2437 9168 2468
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 11756 2468 13277 2496
rect 11756 2456 11762 2468
rect 13265 2465 13277 2468
rect 13311 2465 13323 2499
rect 14550 2496 14556 2508
rect 13265 2459 13323 2465
rect 13832 2468 14556 2496
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 10594 2428 10600 2440
rect 9364 2400 10600 2428
rect 9364 2388 9370 2400
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11020 2400 11253 2428
rect 11020 2388 11026 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 12802 2388 12808 2440
rect 12860 2388 12866 2440
rect 13078 2388 13084 2440
rect 13136 2388 13142 2440
rect 13832 2437 13860 2468
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 13817 2431 13875 2437
rect 13817 2397 13829 2431
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14185 2431 14243 2437
rect 14185 2428 14197 2431
rect 13964 2400 14197 2428
rect 13964 2388 13970 2400
rect 14185 2397 14197 2400
rect 14231 2397 14243 2431
rect 14185 2391 14243 2397
rect 2041 2363 2099 2369
rect 2041 2360 2053 2363
rect 1596 2332 2053 2360
rect 1489 2323 1547 2329
rect 2041 2329 2053 2332
rect 2087 2329 2099 2363
rect 2041 2323 2099 2329
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 9766 2360 9772 2372
rect 8711 2332 9772 2360
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 9766 2320 9772 2332
rect 9824 2320 9830 2372
rect 14553 2363 14611 2369
rect 14553 2329 14565 2363
rect 14599 2360 14611 2363
rect 15470 2360 15476 2372
rect 14599 2332 15476 2360
rect 14599 2329 14611 2332
rect 14553 2323 14611 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 6454 2252 6460 2304
rect 6512 2252 6518 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 1104 2202 14904 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 14904 2202
rect 1104 2128 14904 2150
<< via1 >>
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 14214 15750 14266 15802
rect 14278 15750 14330 15802
rect 14342 15750 14394 15802
rect 14406 15750 14458 15802
rect 14470 15750 14522 15802
rect 940 15648 992 15700
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 10416 15648 10468 15700
rect 20 15444 72 15496
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 9036 15444 9088 15496
rect 11612 15444 11664 15496
rect 13544 15444 13596 15496
rect 15476 15444 15528 15496
rect 5724 15376 5776 15428
rect 7656 15376 7708 15428
rect 2136 15351 2188 15360
rect 2136 15317 2145 15351
rect 2145 15317 2179 15351
rect 2179 15317 2188 15351
rect 2136 15308 2188 15317
rect 2872 15351 2924 15360
rect 2872 15317 2881 15351
rect 2881 15317 2915 15351
rect 2915 15317 2924 15351
rect 2872 15308 2924 15317
rect 4804 15351 4856 15360
rect 4804 15317 4813 15351
rect 4813 15317 4847 15351
rect 4847 15317 4856 15351
rect 4804 15308 4856 15317
rect 8760 15308 8812 15360
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 13728 15351 13780 15360
rect 13728 15317 13737 15351
rect 13737 15317 13771 15351
rect 13771 15317 13780 15351
rect 13728 15308 13780 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 14832 15104 14884 15156
rect 13820 14968 13872 15020
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 14214 14662 14266 14714
rect 14278 14662 14330 14714
rect 14342 14662 14394 14714
rect 14406 14662 14458 14714
rect 14470 14662 14522 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 7932 13880 7984 13932
rect 13912 13880 13964 13932
rect 6552 13812 6604 13864
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 14832 13812 14884 13864
rect 8208 13744 8260 13796
rect 8484 13676 8536 13728
rect 9588 13676 9640 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 14214 13574 14266 13626
rect 14278 13574 14330 13626
rect 14342 13574 14394 13626
rect 14406 13574 14458 13626
rect 14470 13574 14522 13626
rect 4804 13472 4856 13524
rect 5448 13472 5500 13524
rect 6552 13472 6604 13524
rect 9496 13472 9548 13524
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 6000 13336 6052 13388
rect 5356 13268 5408 13320
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 6736 13268 6788 13320
rect 8484 13404 8536 13456
rect 7748 13336 7800 13388
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 9128 13379 9180 13388
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 9588 13336 9640 13388
rect 10416 13404 10468 13456
rect 9220 13311 9272 13320
rect 7932 13200 7984 13252
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9864 13311 9916 13320
rect 9220 13268 9272 13277
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10416 13268 10468 13320
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 7840 13132 7892 13184
rect 10048 13200 10100 13252
rect 9680 13132 9732 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 4712 12928 4764 12980
rect 5264 12903 5316 12912
rect 5264 12869 5273 12903
rect 5273 12869 5307 12903
rect 5307 12869 5316 12903
rect 5264 12860 5316 12869
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 4712 12792 4764 12844
rect 5356 12792 5408 12844
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 8024 12928 8076 12980
rect 8300 12928 8352 12980
rect 9128 12928 9180 12980
rect 9680 12928 9732 12980
rect 10140 12928 10192 12980
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 9864 12860 9916 12912
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 8024 12792 8076 12844
rect 10968 12792 11020 12844
rect 8392 12656 8444 12708
rect 11336 12656 11388 12708
rect 13728 12792 13780 12844
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 14214 12486 14266 12538
rect 14278 12486 14330 12538
rect 14342 12486 14394 12538
rect 14406 12486 14458 12538
rect 14470 12486 14522 12538
rect 5908 12248 5960 12300
rect 4712 12180 4764 12232
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 9956 12180 10008 12232
rect 6368 12112 6420 12164
rect 8760 12112 8812 12164
rect 13912 12112 13964 12164
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 7196 12044 7248 12096
rect 11060 12044 11112 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 3884 11840 3936 11892
rect 4620 11840 4672 11892
rect 6092 11840 6144 11892
rect 940 11704 992 11756
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 5448 11772 5500 11824
rect 8300 11840 8352 11892
rect 8760 11840 8812 11892
rect 4712 11704 4764 11756
rect 4804 11704 4856 11756
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 6276 11772 6328 11824
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 7380 11704 7432 11756
rect 4068 11568 4120 11620
rect 6552 11679 6604 11688
rect 6552 11645 6561 11679
rect 6561 11645 6595 11679
rect 6595 11645 6604 11679
rect 6552 11636 6604 11645
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 9956 11815 10008 11824
rect 9956 11781 9965 11815
rect 9965 11781 9999 11815
rect 9999 11781 10008 11815
rect 9956 11772 10008 11781
rect 11060 11883 11112 11892
rect 11060 11849 11069 11883
rect 11069 11849 11103 11883
rect 11103 11849 11112 11883
rect 11060 11840 11112 11849
rect 7196 11500 7248 11552
rect 7564 11543 7616 11552
rect 7564 11509 7573 11543
rect 7573 11509 7607 11543
rect 7607 11509 7616 11543
rect 7564 11500 7616 11509
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 8116 11636 8168 11688
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 9772 11747 9824 11756
rect 9772 11713 9779 11747
rect 9779 11713 9824 11747
rect 8852 11636 8904 11688
rect 7932 11568 7984 11620
rect 9220 11679 9272 11688
rect 9220 11645 9229 11679
rect 9229 11645 9263 11679
rect 9263 11645 9272 11679
rect 9220 11636 9272 11645
rect 9772 11704 9824 11713
rect 10048 11747 10100 11756
rect 10048 11713 10062 11747
rect 10062 11713 10096 11747
rect 10096 11713 10100 11747
rect 10048 11704 10100 11713
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 9864 11636 9916 11688
rect 13820 11568 13872 11620
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 14214 11398 14266 11450
rect 14278 11398 14330 11450
rect 14342 11398 14394 11450
rect 14406 11398 14458 11450
rect 14470 11398 14522 11450
rect 5632 11296 5684 11348
rect 6092 11296 6144 11348
rect 6552 11296 6604 11348
rect 7288 11296 7340 11348
rect 3884 11092 3936 11144
rect 4160 11160 4212 11212
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 6368 11024 6420 11076
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8024 11092 8076 11144
rect 9220 11296 9272 11348
rect 10784 11296 10836 11348
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 9680 11228 9732 11280
rect 8300 11160 8352 11212
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 9588 11135 9640 11144
rect 9588 11101 9597 11135
rect 9597 11101 9631 11135
rect 9631 11101 9640 11135
rect 9588 11092 9640 11101
rect 10600 11092 10652 11144
rect 8576 11024 8628 11076
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 11152 11092 11204 11101
rect 11244 11092 11296 11144
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 6552 10956 6604 11008
rect 11704 11024 11756 11076
rect 14924 11024 14976 11076
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 4804 10752 4856 10804
rect 8208 10752 8260 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 7288 10684 7340 10736
rect 7840 10727 7892 10736
rect 7840 10693 7849 10727
rect 7849 10693 7883 10727
rect 7883 10693 7892 10727
rect 7840 10684 7892 10693
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 3884 10548 3936 10600
rect 2228 10480 2280 10532
rect 6920 10616 6972 10668
rect 10968 10616 11020 10668
rect 11612 10616 11664 10668
rect 4804 10480 4856 10532
rect 9312 10480 9364 10532
rect 6276 10412 6328 10464
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 8300 10412 8352 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 14214 10310 14266 10362
rect 14278 10310 14330 10362
rect 14342 10310 14394 10362
rect 14406 10310 14458 10362
rect 14470 10310 14522 10362
rect 8300 10208 8352 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 9496 10208 9548 10260
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 5448 10140 5500 10192
rect 7472 10140 7524 10192
rect 4804 10072 4856 10124
rect 5264 10004 5316 10056
rect 4344 9979 4396 9988
rect 4344 9945 4353 9979
rect 4353 9945 4387 9979
rect 4387 9945 4396 9979
rect 4344 9936 4396 9945
rect 6092 10004 6144 10056
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 10232 10208 10284 10260
rect 10968 10208 11020 10260
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 6644 10004 6696 10056
rect 5816 9936 5868 9988
rect 6276 9936 6328 9988
rect 6368 9936 6420 9988
rect 6920 10004 6972 10056
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 7288 10047 7340 10056
rect 7288 10013 7300 10047
rect 7300 10013 7334 10047
rect 7334 10013 7340 10047
rect 7288 10004 7340 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 9588 10072 9640 10124
rect 9864 10004 9916 10056
rect 7932 9936 7984 9988
rect 8760 9936 8812 9988
rect 4620 9868 4672 9920
rect 6828 9868 6880 9920
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 10232 9936 10284 9988
rect 10048 9868 10100 9920
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 11336 10004 11388 10056
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 11980 9936 12032 9988
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 4068 9664 4120 9716
rect 4344 9664 4396 9716
rect 5816 9664 5868 9716
rect 6368 9596 6420 9648
rect 6736 9664 6788 9716
rect 8024 9664 8076 9716
rect 9220 9707 9272 9716
rect 9220 9673 9229 9707
rect 9229 9673 9263 9707
rect 9263 9673 9272 9707
rect 9220 9664 9272 9673
rect 9588 9664 9640 9716
rect 4712 9528 4764 9580
rect 6092 9528 6144 9580
rect 6828 9596 6880 9648
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 4620 9460 4672 9512
rect 5172 9460 5224 9512
rect 7012 9460 7064 9512
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 7472 9528 7524 9537
rect 7932 9528 7984 9580
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 9680 9596 9732 9648
rect 9956 9639 10008 9648
rect 9956 9605 9965 9639
rect 9965 9605 9999 9639
rect 9999 9605 10008 9639
rect 9956 9596 10008 9605
rect 10232 9634 10284 9686
rect 8116 9392 8168 9444
rect 9312 9460 9364 9512
rect 10048 9528 10100 9580
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 10968 9528 11020 9580
rect 11060 9528 11112 9580
rect 11244 9528 11296 9580
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 10784 9460 10836 9512
rect 12808 9460 12860 9512
rect 3700 9324 3752 9376
rect 4344 9324 4396 9376
rect 4804 9324 4856 9376
rect 7748 9324 7800 9376
rect 8208 9324 8260 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 14214 9222 14266 9274
rect 14278 9222 14330 9274
rect 14342 9222 14394 9274
rect 14406 9222 14458 9274
rect 14470 9222 14522 9274
rect 6920 9120 6972 9172
rect 7196 9120 7248 9172
rect 7656 9120 7708 9172
rect 10048 9120 10100 9172
rect 10232 9120 10284 9172
rect 10784 9120 10836 9172
rect 10876 9163 10928 9172
rect 10876 9129 10885 9163
rect 10885 9129 10919 9163
rect 10919 9129 10928 9163
rect 10876 9120 10928 9129
rect 4344 9052 4396 9104
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 5724 9052 5776 9104
rect 6828 9052 6880 9104
rect 8208 9052 8260 9104
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 4620 8959 4672 8968
rect 4620 8925 4627 8959
rect 4627 8925 4672 8959
rect 4620 8916 4672 8925
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5172 8916 5224 8968
rect 5448 8916 5500 8968
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 6552 8916 6604 8968
rect 940 8848 992 8900
rect 5356 8848 5408 8900
rect 6828 8916 6880 8968
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 5448 8780 5500 8832
rect 5816 8823 5868 8832
rect 5816 8789 5825 8823
rect 5825 8789 5859 8823
rect 5859 8789 5868 8823
rect 5816 8780 5868 8789
rect 6644 8780 6696 8832
rect 6736 8823 6788 8832
rect 6736 8789 6745 8823
rect 6745 8789 6779 8823
rect 6779 8789 6788 8823
rect 6736 8780 6788 8789
rect 6920 8780 6972 8832
rect 7748 8780 7800 8832
rect 9864 8916 9916 8968
rect 9772 8848 9824 8900
rect 10324 8823 10376 8832
rect 10324 8789 10333 8823
rect 10333 8789 10367 8823
rect 10367 8789 10376 8823
rect 10324 8780 10376 8789
rect 11520 9163 11572 9172
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 11888 8984 11940 9036
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 13268 8916 13320 8968
rect 11796 8891 11848 8900
rect 11796 8857 11805 8891
rect 11805 8857 11839 8891
rect 11839 8857 11848 8891
rect 11796 8848 11848 8857
rect 10968 8780 11020 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 12164 8823 12216 8832
rect 12164 8789 12173 8823
rect 12173 8789 12207 8823
rect 12207 8789 12216 8823
rect 12164 8780 12216 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4068 8576 4120 8628
rect 4436 8576 4488 8628
rect 3792 8508 3844 8560
rect 4344 8508 4396 8560
rect 4804 8440 4856 8492
rect 5540 8576 5592 8628
rect 5816 8576 5868 8628
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 7380 8576 7432 8628
rect 5356 8508 5408 8560
rect 5448 8508 5500 8560
rect 6552 8508 6604 8560
rect 7656 8576 7708 8628
rect 9588 8576 9640 8628
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 7472 8440 7524 8492
rect 11152 8576 11204 8628
rect 11796 8576 11848 8628
rect 11888 8576 11940 8628
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 9404 8440 9456 8492
rect 9772 8440 9824 8492
rect 9956 8440 10008 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 9680 8372 9732 8424
rect 3424 8279 3476 8288
rect 3424 8245 3433 8279
rect 3433 8245 3467 8279
rect 3467 8245 3476 8279
rect 3424 8236 3476 8245
rect 3884 8236 3936 8288
rect 6552 8304 6604 8356
rect 9496 8304 9548 8356
rect 9956 8347 10008 8356
rect 9956 8313 9965 8347
rect 9965 8313 9999 8347
rect 9999 8313 10008 8347
rect 9956 8304 10008 8313
rect 10692 8440 10744 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 12164 8508 12216 8560
rect 12808 8440 12860 8492
rect 14464 8551 14516 8560
rect 14464 8517 14473 8551
rect 14473 8517 14507 8551
rect 14507 8517 14516 8551
rect 14464 8508 14516 8517
rect 5172 8236 5224 8288
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 6828 8236 6880 8288
rect 10692 8304 10744 8356
rect 11244 8304 11296 8356
rect 11336 8304 11388 8356
rect 11612 8304 11664 8356
rect 10968 8236 11020 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 14214 8134 14266 8186
rect 14278 8134 14330 8186
rect 14342 8134 14394 8186
rect 14406 8134 14458 8186
rect 14470 8134 14522 8186
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 8392 8032 8444 8084
rect 9128 8032 9180 8084
rect 5172 7964 5224 8016
rect 3424 7896 3476 7948
rect 2872 7828 2924 7880
rect 3884 7871 3936 7880
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 5264 7896 5316 7948
rect 7472 7896 7524 7948
rect 7840 7896 7892 7948
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 8760 7896 8812 7948
rect 4068 7828 4120 7880
rect 5356 7828 5408 7880
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 6828 7828 6880 7880
rect 4436 7760 4488 7812
rect 7196 7828 7248 7880
rect 3516 7692 3568 7744
rect 4620 7692 4672 7744
rect 4804 7692 4856 7744
rect 5356 7692 5408 7744
rect 6644 7692 6696 7744
rect 6920 7692 6972 7744
rect 8852 7828 8904 7880
rect 9312 7828 9364 7880
rect 10508 7896 10560 7948
rect 12808 7896 12860 7948
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 10048 7828 10100 7880
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 8208 7692 8260 7744
rect 9036 7692 9088 7744
rect 10600 7692 10652 7744
rect 11796 7692 11848 7744
rect 13268 7692 13320 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 3976 7420 4028 7472
rect 5264 7420 5316 7472
rect 5448 7420 5500 7472
rect 6460 7463 6512 7472
rect 6460 7429 6469 7463
rect 6469 7429 6503 7463
rect 6503 7429 6512 7463
rect 6460 7420 6512 7429
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 3424 7352 3476 7404
rect 3700 7352 3752 7404
rect 3884 7352 3936 7404
rect 4620 7352 4672 7404
rect 6552 7352 6604 7404
rect 3608 7216 3660 7268
rect 4712 7216 4764 7268
rect 7840 7488 7892 7540
rect 7932 7488 7984 7540
rect 8760 7531 8812 7540
rect 8760 7497 8769 7531
rect 8769 7497 8803 7531
rect 8803 7497 8812 7531
rect 8760 7488 8812 7497
rect 9128 7488 9180 7540
rect 10140 7488 10192 7540
rect 9404 7420 9456 7472
rect 8852 7352 8904 7404
rect 9036 7352 9088 7404
rect 11244 7420 11296 7472
rect 11428 7420 11480 7472
rect 10416 7352 10468 7404
rect 10784 7352 10836 7404
rect 10876 7352 10928 7404
rect 11152 7352 11204 7404
rect 11980 7352 12032 7404
rect 10232 7284 10284 7336
rect 11520 7284 11572 7336
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 5264 7148 5316 7200
rect 6644 7148 6696 7200
rect 6828 7148 6880 7200
rect 7012 7148 7064 7200
rect 8392 7148 8444 7200
rect 9680 7148 9732 7200
rect 10692 7148 10744 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 14214 7046 14266 7098
rect 14278 7046 14330 7098
rect 14342 7046 14394 7098
rect 14406 7046 14458 7098
rect 14470 7046 14522 7098
rect 2872 6740 2924 6792
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 3240 6740 3292 6792
rect 4620 6944 4672 6996
rect 3608 6876 3660 6928
rect 3792 6851 3844 6860
rect 3792 6817 3801 6851
rect 3801 6817 3835 6851
rect 3835 6817 3844 6851
rect 3792 6808 3844 6817
rect 3516 6740 3568 6792
rect 4068 6740 4120 6792
rect 4804 6876 4856 6928
rect 5724 6944 5776 6996
rect 4252 6808 4304 6860
rect 4712 6808 4764 6860
rect 8944 6944 8996 6996
rect 10876 6944 10928 6996
rect 11704 6944 11756 6996
rect 6828 6876 6880 6928
rect 5908 6808 5960 6860
rect 8576 6808 8628 6860
rect 10692 6876 10744 6928
rect 4528 6740 4580 6792
rect 4896 6740 4948 6792
rect 5448 6672 5500 6724
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6644 6740 6696 6792
rect 8484 6740 8536 6792
rect 5724 6604 5776 6656
rect 6460 6672 6512 6724
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6000 6604 6052 6613
rect 6368 6604 6420 6656
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 9220 6604 9272 6656
rect 9680 6740 9732 6792
rect 9680 6604 9732 6656
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 9864 6604 9916 6656
rect 10140 6740 10192 6792
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 10416 6604 10468 6656
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 10876 6740 10928 6749
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 10600 6715 10652 6724
rect 10600 6681 10609 6715
rect 10609 6681 10643 6715
rect 10643 6681 10652 6715
rect 10600 6672 10652 6681
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 11612 6740 11664 6792
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 3884 6400 3936 6452
rect 4252 6400 4304 6452
rect 3976 6332 4028 6384
rect 4528 6332 4580 6384
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 5540 6400 5592 6452
rect 6000 6400 6052 6452
rect 6644 6400 6696 6452
rect 7012 6400 7064 6452
rect 7104 6400 7156 6452
rect 10692 6400 10744 6452
rect 10968 6400 11020 6452
rect 11152 6400 11204 6452
rect 3424 6264 3476 6316
rect 3332 6196 3384 6248
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 3240 6060 3292 6112
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 3792 6060 3844 6112
rect 6920 6264 6972 6316
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 6552 6128 6604 6180
rect 7932 6196 7984 6248
rect 8760 6264 8812 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 9864 6332 9916 6384
rect 12624 6400 12676 6452
rect 13360 6400 13412 6452
rect 9036 6264 9088 6316
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 4712 6060 4764 6112
rect 8208 6060 8260 6112
rect 8852 6128 8904 6180
rect 10508 6264 10560 6316
rect 10784 6264 10836 6316
rect 11888 6264 11940 6316
rect 9404 6196 9456 6248
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 14924 6264 14976 6316
rect 9588 6060 9640 6112
rect 12440 6128 12492 6180
rect 11060 6060 11112 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 14214 5958 14266 6010
rect 14278 5958 14330 6010
rect 14342 5958 14394 6010
rect 14406 5958 14458 6010
rect 14470 5958 14522 6010
rect 3332 5856 3384 5908
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 7012 5899 7064 5908
rect 7012 5865 7021 5899
rect 7021 5865 7055 5899
rect 7055 5865 7064 5899
rect 7012 5856 7064 5865
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 9036 5856 9088 5908
rect 9588 5856 9640 5908
rect 10600 5856 10652 5908
rect 12440 5899 12492 5908
rect 12440 5865 12449 5899
rect 12449 5865 12483 5899
rect 12483 5865 12492 5899
rect 12440 5856 12492 5865
rect 2136 5720 2188 5772
rect 4804 5720 4856 5772
rect 3424 5652 3476 5704
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 3148 5584 3200 5636
rect 7840 5652 7892 5704
rect 10324 5788 10376 5840
rect 12808 5788 12860 5840
rect 9220 5720 9272 5772
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 8024 5584 8076 5636
rect 8392 5627 8444 5636
rect 8392 5593 8401 5627
rect 8401 5593 8435 5627
rect 8435 5593 8444 5627
rect 8392 5584 8444 5593
rect 13820 5720 13872 5772
rect 11336 5695 11388 5704
rect 11336 5661 11355 5695
rect 11355 5661 11388 5695
rect 11336 5652 11388 5661
rect 11796 5652 11848 5704
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 10600 5584 10652 5636
rect 11520 5627 11572 5636
rect 11520 5593 11529 5627
rect 11529 5593 11563 5627
rect 11563 5593 11572 5627
rect 11520 5584 11572 5593
rect 12440 5584 12492 5636
rect 9404 5516 9456 5568
rect 11060 5516 11112 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5816 5312 5868 5364
rect 5356 5287 5408 5296
rect 5356 5253 5365 5287
rect 5365 5253 5399 5287
rect 5399 5253 5408 5287
rect 5356 5244 5408 5253
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 5264 5176 5316 5228
rect 5448 5176 5500 5228
rect 5724 5176 5776 5228
rect 6828 5312 6880 5364
rect 5356 5040 5408 5092
rect 4620 4972 4672 5024
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 7012 5176 7064 5228
rect 8208 5244 8260 5296
rect 8392 5244 8444 5296
rect 8116 5176 8168 5228
rect 9956 5176 10008 5228
rect 10232 5176 10284 5228
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 10600 5176 10652 5228
rect 10692 5176 10744 5228
rect 8484 5108 8536 5160
rect 9404 5108 9456 5160
rect 10048 5151 10100 5160
rect 10048 5117 10057 5151
rect 10057 5117 10091 5151
rect 10091 5117 10100 5151
rect 10048 5108 10100 5117
rect 10324 5151 10376 5160
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 11152 5312 11204 5364
rect 12440 5312 12492 5364
rect 13360 5355 13412 5364
rect 13360 5321 13369 5355
rect 13369 5321 13403 5355
rect 13403 5321 13412 5355
rect 13360 5312 13412 5321
rect 11244 5287 11296 5296
rect 11244 5253 11253 5287
rect 11253 5253 11287 5287
rect 11287 5253 11296 5287
rect 11244 5244 11296 5253
rect 12532 5176 12584 5228
rect 11152 5151 11204 5160
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 8024 5015 8076 5024
rect 8024 4981 8033 5015
rect 8033 4981 8067 5015
rect 8067 4981 8076 5015
rect 8024 4972 8076 4981
rect 9128 4972 9180 5024
rect 9588 4972 9640 5024
rect 10324 4972 10376 5024
rect 11612 4972 11664 5024
rect 13268 5040 13320 5092
rect 13176 5015 13228 5024
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 14214 4870 14266 4922
rect 14278 4870 14330 4922
rect 14342 4870 14394 4922
rect 14406 4870 14458 4922
rect 14470 4870 14522 4922
rect 6368 4768 6420 4820
rect 7656 4768 7708 4820
rect 7932 4768 7984 4820
rect 8024 4768 8076 4820
rect 5816 4700 5868 4752
rect 6828 4700 6880 4752
rect 7748 4700 7800 4752
rect 940 4564 992 4616
rect 4804 4564 4856 4616
rect 5356 4564 5408 4616
rect 8576 4632 8628 4684
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 6828 4564 6880 4616
rect 7748 4564 7800 4616
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 10692 4700 10744 4752
rect 11520 4768 11572 4820
rect 12440 4768 12492 4820
rect 13820 4768 13872 4820
rect 11428 4700 11480 4752
rect 10048 4564 10100 4616
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 11704 4564 11756 4616
rect 4804 4428 4856 4480
rect 5540 4428 5592 4480
rect 6368 4471 6420 4480
rect 6368 4437 6377 4471
rect 6377 4437 6411 4471
rect 6411 4437 6420 4471
rect 6368 4428 6420 4437
rect 6460 4428 6512 4480
rect 6920 4428 6972 4480
rect 7012 4428 7064 4480
rect 9036 4428 9088 4480
rect 9220 4428 9272 4480
rect 10508 4428 10560 4480
rect 14924 4428 14976 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5540 4224 5592 4276
rect 8208 4224 8260 4276
rect 8300 4224 8352 4276
rect 9036 4224 9088 4276
rect 13912 4224 13964 4276
rect 4620 4088 4672 4140
rect 4804 4131 4856 4140
rect 4804 4097 4814 4131
rect 4814 4097 4848 4131
rect 4848 4097 4856 4131
rect 4804 4088 4856 4097
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 5356 4088 5408 4140
rect 5816 4020 5868 4072
rect 5448 3884 5500 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 7748 3884 7800 3936
rect 8116 3952 8168 4004
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 9496 4088 9548 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 10048 4088 10100 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 10324 4156 10376 4208
rect 11520 4156 11572 4208
rect 12072 4088 12124 4140
rect 8392 4020 8444 4029
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 8484 3952 8536 4004
rect 9312 3884 9364 3936
rect 9680 3884 9732 3936
rect 10784 3884 10836 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 14214 3782 14266 3834
rect 14278 3782 14330 3834
rect 14342 3782 14394 3834
rect 14406 3782 14458 3834
rect 14470 3782 14522 3834
rect 4988 3680 5040 3732
rect 5264 3612 5316 3664
rect 6460 3612 6512 3664
rect 6644 3612 6696 3664
rect 6920 3612 6972 3664
rect 7840 3723 7892 3732
rect 7840 3689 7849 3723
rect 7849 3689 7883 3723
rect 7883 3689 7892 3723
rect 7840 3680 7892 3689
rect 9864 3680 9916 3732
rect 10140 3680 10192 3732
rect 11796 3680 11848 3732
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 7656 3544 7708 3596
rect 10324 3612 10376 3664
rect 8668 3476 8720 3528
rect 9680 3476 9732 3528
rect 5356 3408 5408 3460
rect 5540 3408 5592 3460
rect 6828 3408 6880 3460
rect 9588 3451 9640 3460
rect 9588 3417 9597 3451
rect 9597 3417 9631 3451
rect 9631 3417 9640 3451
rect 9588 3408 9640 3417
rect 4804 3340 4856 3392
rect 8944 3340 8996 3392
rect 12072 3655 12124 3664
rect 12072 3621 12081 3655
rect 12081 3621 12115 3655
rect 12115 3621 12124 3655
rect 12072 3612 12124 3621
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 10508 3451 10560 3460
rect 10508 3417 10517 3451
rect 10517 3417 10551 3451
rect 10551 3417 10560 3451
rect 10508 3408 10560 3417
rect 10416 3340 10468 3392
rect 11704 3451 11756 3460
rect 11704 3417 11713 3451
rect 11713 3417 11747 3451
rect 11747 3417 11756 3451
rect 11704 3408 11756 3417
rect 12532 3340 12584 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5264 3136 5316 3188
rect 3976 3000 4028 3052
rect 4804 3000 4856 3052
rect 5356 3000 5408 3052
rect 5632 3068 5684 3120
rect 6092 3136 6144 3188
rect 6368 3000 6420 3052
rect 6460 3000 6512 3052
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 7656 3000 7708 3052
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8576 3068 8628 3120
rect 6828 2932 6880 2941
rect 7748 2864 7800 2916
rect 9588 3136 9640 3188
rect 9956 3136 10008 3188
rect 10324 3136 10376 3188
rect 8944 3111 8996 3120
rect 8944 3077 8953 3111
rect 8953 3077 8987 3111
rect 8987 3077 8996 3111
rect 8944 3068 8996 3077
rect 10048 3111 10100 3120
rect 10048 3077 10057 3111
rect 10057 3077 10091 3111
rect 10091 3077 10100 3111
rect 10048 3068 10100 3077
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 10600 3043 10652 3052
rect 10600 3009 10617 3043
rect 10617 3009 10651 3043
rect 10651 3009 10652 3043
rect 10600 3000 10652 3009
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 13176 3068 13228 3120
rect 12532 3000 12584 3052
rect 8668 2839 8720 2848
rect 8668 2805 8677 2839
rect 8677 2805 8711 2839
rect 8711 2805 8720 2839
rect 8668 2796 8720 2805
rect 10784 2796 10836 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 14214 2694 14266 2746
rect 14278 2694 14330 2746
rect 14342 2694 14394 2746
rect 14406 2694 14458 2746
rect 14470 2694 14522 2746
rect 2228 2592 2280 2644
rect 2872 2592 2924 2644
rect 4068 2592 4120 2644
rect 6184 2592 6236 2644
rect 7840 2592 7892 2644
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 7748 2567 7800 2576
rect 7748 2533 7757 2567
rect 7757 2533 7791 2567
rect 7791 2533 7800 2567
rect 7748 2524 7800 2533
rect 8668 2456 8720 2508
rect 20 2388 72 2440
rect 940 2320 992 2372
rect 1952 2388 2004 2440
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 10784 2456 10836 2508
rect 11704 2456 11756 2508
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 10600 2388 10652 2440
rect 10968 2388 11020 2440
rect 12808 2431 12860 2440
rect 12808 2397 12817 2431
rect 12817 2397 12851 2431
rect 12851 2397 12860 2431
rect 12808 2388 12860 2397
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 14556 2456 14608 2508
rect 13912 2388 13964 2440
rect 9772 2320 9824 2372
rect 15476 2320 15528 2372
rect 6460 2295 6512 2304
rect 6460 2261 6469 2295
rect 6469 2261 6503 2295
rect 6503 2261 6512 2295
rect 6460 2252 6512 2261
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 18 17433 74 18233
rect 2594 17433 2650 18233
rect 4526 17433 4582 18233
rect 7102 17433 7158 18233
rect 9034 17433 9090 18233
rect 11610 17433 11666 18233
rect 13542 17433 13598 18233
rect 15474 17433 15530 18233
rect 32 15502 60 17433
rect 2608 16574 2636 17433
rect 4540 16574 4568 17433
rect 7116 16574 7144 17433
rect 2608 16546 2728 16574
rect 4540 16546 4660 16574
rect 7116 16546 7328 16574
rect 938 16416 994 16425
rect 938 16351 994 16360
rect 952 15706 980 16351
rect 940 15700 992 15706
rect 940 15642 992 15648
rect 2700 15502 2728 16546
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15502 4660 16546
rect 7300 15706 7328 16546
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 9048 15502 9076 17433
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 20 15496 72 15502
rect 20 15438 72 15444
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 938 8936 994 8945
rect 938 8871 940 8880
rect 992 8871 994 8880
rect 940 8842 992 8848
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6905 1532 7346
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 2148 5778 2176 15302
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4185 980 4558
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 2240 2650 2268 10474
rect 2884 7886 2912 15302
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4816 13530 4844 15302
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4724 12986 4752 13126
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 11898 4660 12786
rect 4724 12238 4752 12786
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 3896 11762 3924 11834
rect 4724 11762 4752 12174
rect 4816 11762 4844 13466
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5276 12918 5304 13330
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5368 12850 5396 13262
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5460 11830 5488 13466
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 3896 11150 3924 11698
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4080 11234 4108 11562
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4080 11218 4200 11234
rect 4080 11212 4212 11218
rect 4080 11206 4160 11212
rect 4160 11154 4212 11160
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3896 10606 3924 11086
rect 4172 10674 4200 11154
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 10810 4844 11086
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3896 9518 3924 10542
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4816 10130 4844 10474
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 4080 9722 4108 9998
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4356 9722 4384 9930
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 4356 9382 4384 9658
rect 4632 9518 4660 9862
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7954 3464 8230
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2884 6798 2912 7822
rect 3436 7410 3464 7890
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3528 6798 3556 7686
rect 3712 7410 3740 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 4080 8634 4108 8871
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4356 8566 4384 9046
rect 4632 8974 4660 9454
rect 4724 8974 4752 9522
rect 5172 9512 5224 9518
rect 5276 9500 5304 9998
rect 5224 9472 5304 9500
rect 5172 9454 5224 9460
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4448 8634 4476 8910
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3620 6934 3648 7210
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3804 6866 3832 8502
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 7886 3924 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3896 7410 3924 7822
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 2650 2912 6054
rect 3160 5642 3188 6734
rect 3252 6118 3280 6734
rect 3424 6316 3476 6322
rect 3804 6304 3832 6802
rect 3896 6458 3924 7346
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3988 6390 4016 7414
rect 4080 6882 4108 7822
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4448 7206 4476 7754
rect 4632 7750 4660 8910
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4724 7426 4752 8910
rect 4816 8498 4844 9318
rect 5184 8974 5212 9454
rect 5368 9042 5396 11698
rect 5460 10198 5488 11766
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11354 5672 11698
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5460 8974 5488 10134
rect 5736 9110 5764 15370
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 6564 13530 6592 13806
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5920 11762 5948 12242
rect 6012 11762 6040 13330
rect 6564 13326 6592 13466
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6104 11898 6132 12174
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5814 10024 5870 10033
rect 5814 9959 5816 9968
rect 5868 9959 5870 9968
rect 5816 9930 5868 9936
rect 5828 9722 5856 9930
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5172 8968 5224 8974
rect 5448 8968 5500 8974
rect 5224 8928 5304 8956
rect 5172 8910 5224 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4816 7750 4844 8434
rect 5276 8378 5304 8928
rect 5448 8910 5500 8916
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 8566 5396 8842
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8566 5488 8774
rect 5552 8634 5580 8910
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5276 8350 5396 8378
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5184 8022 5212 8230
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5184 7834 5212 7958
rect 5276 7954 5304 8230
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5368 7886 5396 8350
rect 5356 7880 5408 7886
rect 5184 7806 5304 7834
rect 5356 7822 5408 7828
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7478 5304 7806
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5264 7472 5316 7478
rect 4620 7404 4672 7410
rect 4724 7398 4936 7426
rect 5264 7414 5316 7420
rect 4620 7346 4672 7352
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 7002 4660 7346
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4080 6866 4292 6882
rect 4724 6866 4752 7210
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4080 6860 4304 6866
rect 4080 6854 4252 6860
rect 4252 6802 4304 6808
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3476 6276 3832 6304
rect 3424 6258 3476 6264
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3344 5914 3372 6190
rect 3804 6118 3832 6276
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3436 5710 3464 6054
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 3058 4016 5510
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4080 2650 4108 6734
rect 4264 6458 4292 6802
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4540 6390 4568 6734
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4724 6118 4752 6802
rect 4816 6458 4844 6870
rect 4908 6798 4936 7398
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4816 5234 4844 5714
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5276 5234 5304 7142
rect 5368 6610 5396 7686
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5460 6730 5488 7414
rect 5644 7018 5672 8910
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8634 5856 8774
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5920 7018 5948 11698
rect 6104 11354 6132 11834
rect 6288 11830 6316 12038
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6380 11082 6408 12106
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6564 11354 6592 11630
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6104 9586 6132 9998
rect 6288 9994 6316 10406
rect 6564 10062 6592 10950
rect 6748 10130 6776 13262
rect 7392 12986 7420 13806
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5552 6990 5672 7018
rect 5736 7002 5948 7018
rect 5724 6996 5948 7002
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5368 6582 5488 6610
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5368 5302 5396 5850
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4146 4660 4966
rect 4816 4622 4844 5170
rect 5368 5098 5396 5238
rect 5460 5234 5488 6582
rect 5552 6458 5580 6990
rect 5776 6990 5948 6996
rect 5724 6938 5776 6944
rect 5920 6866 5948 6990
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6662 5764 6734
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6012 6458 6040 6598
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5552 5114 5580 6394
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5736 5137 5764 5170
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5460 5086 5580 5114
rect 5722 5128 5778 5137
rect 5368 4622 5396 5034
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4146 4844 4422
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5460 4162 5488 5086
rect 5722 5063 5778 5072
rect 5828 4758 5856 5306
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4282 5580 4422
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5368 4146 5488 4162
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5356 4140 5488 4146
rect 5408 4134 5488 4140
rect 5356 4082 5408 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5000 3738 5028 4082
rect 5828 4078 5856 4694
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5906 4040 5962 4049
rect 5906 3975 5962 3984
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4816 3058 4844 3334
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5276 3194 5304 3606
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5368 3058 5396 3402
rect 5460 3210 5488 3878
rect 5552 3466 5580 3878
rect 5920 3602 5948 3975
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5460 3182 5672 3210
rect 6104 3194 6132 3470
rect 5644 3126 5672 3182
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 6288 2774 6316 9930
rect 6380 9654 6408 9930
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6564 8974 6592 9998
rect 6656 9602 6684 9998
rect 6748 9722 6776 10066
rect 6840 9926 6868 11630
rect 7208 11558 7236 12038
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6932 10062 6960 10610
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6828 9648 6880 9654
rect 6656 9596 6828 9602
rect 6656 9590 6880 9596
rect 6656 9574 6868 9590
rect 7024 9518 7052 9998
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7208 9178 7236 11494
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7300 11150 7328 11290
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7300 10062 7328 10678
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6840 8974 6868 9046
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6656 8634 6684 8774
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6564 8362 6592 8502
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 8090 6592 8298
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6472 7478 6500 7822
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6472 6882 6500 7414
rect 6564 7410 6592 8026
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6380 6854 6500 6882
rect 6380 6662 6408 6854
rect 6564 6746 6592 7346
rect 6656 7206 6684 7686
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 6798 6684 7142
rect 6472 6730 6592 6746
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6460 6724 6592 6730
rect 6512 6718 6592 6724
rect 6460 6666 6512 6672
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6564 5710 6592 6122
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4826 6408 5102
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6656 4622 6684 6394
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6380 3534 6408 4422
rect 6472 3670 6500 4422
rect 6656 3670 6684 4558
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6380 3058 6408 3470
rect 6472 3058 6500 3606
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6196 2746 6316 2774
rect 6196 2650 6224 2746
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6748 2446 6776 8774
rect 6840 8401 6868 8910
rect 6932 8838 6960 9114
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 7392 8634 7420 11698
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7484 9586 7512 10134
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7576 8974 7604 11494
rect 7668 9178 7696 15370
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7760 12850 7788 13330
rect 7944 13258 7972 13874
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7852 12594 7880 13126
rect 7944 12850 7972 13194
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8036 12850 8064 12922
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7760 12566 7880 12594
rect 7760 10588 7788 12566
rect 7944 12152 7972 12786
rect 7852 12124 7972 12152
rect 7852 11150 7880 12124
rect 8220 11762 8248 13738
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13462 8524 13670
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8312 12986 8340 13262
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7944 11150 7972 11562
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7852 10742 7880 11086
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7760 10560 7880 10588
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 9382 7788 9862
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7668 8634 7696 9114
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 6826 8392 6882 8401
rect 6826 8327 6882 8336
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 7886 6868 8230
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7206 6868 7822
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6934 6868 7142
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6932 6780 6960 7686
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6840 6752 6960 6780
rect 6840 5370 6868 6752
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6322 6960 6598
rect 7024 6458 7052 7142
rect 7116 6458 7144 8434
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7208 7886 7236 8366
rect 7484 7954 7512 8434
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 5914 7052 6258
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7024 5234 7052 5850
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6840 4622 6868 4694
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6918 4584 6974 4593
rect 6918 4519 6974 4528
rect 6932 4486 6960 4519
rect 7024 4486 7052 4966
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6840 2990 6868 3402
rect 6932 3058 6960 3606
rect 7668 3602 7696 4762
rect 7760 4758 7788 8774
rect 7852 7954 7880 10560
rect 8036 10470 8064 11086
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 7944 9586 7972 9930
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9722 8064 9862
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 8128 9450 8156 11630
rect 8312 11218 8340 11834
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8220 10810 8248 11086
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10266 8340 10406
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9110 8248 9318
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8404 8090 8432 12650
rect 8772 12434 8800 15302
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9140 12986 9168 13330
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9232 12434 9260 13262
rect 8680 12406 8800 12434
rect 9140 12406 9260 12434
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7852 7546 7880 7890
rect 8220 7750 8248 7890
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 7944 7546 7972 7686
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8392 7200 8444 7206
rect 8496 7188 8524 10202
rect 8588 10062 8616 11018
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8680 8945 8708 12406
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8772 11898 8800 12106
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 9140 11762 9168 12406
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 8758 10024 8814 10033
rect 8758 9959 8760 9968
rect 8812 9959 8814 9968
rect 8760 9930 8812 9936
rect 8666 8936 8722 8945
rect 8666 8871 8722 8880
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8772 7546 8800 7890
rect 8864 7886 8892 11630
rect 9232 11354 9260 11630
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9508 11150 9536 13466
rect 9600 13394 9628 13670
rect 10428 13462 10456 15642
rect 11624 15502 11652 17433
rect 13556 15502 13584 17433
rect 14214 15804 14522 15813
rect 14214 15802 14220 15804
rect 14276 15802 14300 15804
rect 14356 15802 14380 15804
rect 14436 15802 14460 15804
rect 14516 15802 14522 15804
rect 14276 15750 14278 15802
rect 14458 15750 14460 15802
rect 14214 15748 14220 15750
rect 14276 15748 14300 15750
rect 14356 15748 14380 15750
rect 14436 15748 14460 15750
rect 14516 15748 14522 15750
rect 14214 15739 14522 15748
rect 14830 15736 14886 15745
rect 14830 15671 14886 15680
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9600 11150 9628 13330
rect 10428 13326 10456 13398
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12986 9720 13126
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9876 12918 9904 13262
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 11830 9996 12174
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10060 11762 10088 13194
rect 10152 12986 10180 13262
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10980 12434 11008 12786
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 10980 12406 11284 12434
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 11898 11100 12038
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 10146 9352 10474
rect 9508 10266 9536 11086
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9324 10130 9628 10146
rect 9324 10124 9640 10130
rect 9324 10118 9588 10124
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9722 9260 9998
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9324 9518 9352 10118
rect 9588 10066 9640 10072
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9508 8945 9536 9522
rect 9494 8936 9550 8945
rect 9494 8871 9550 8880
rect 9600 8634 9628 9658
rect 9692 9654 9720 11222
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9784 9500 9812 11698
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 10266 9904 11630
rect 10796 11354 10824 11698
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 11256 11150 11284 12406
rect 11348 11354 11376 12650
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9692 9472 9812 9500
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9140 8090 9168 8434
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8444 7160 8524 7188
rect 8392 7142 8444 7148
rect 8496 6798 8524 7160
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7944 5914 7972 6190
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7760 3942 7788 4558
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7668 3058 7696 3538
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 7760 2922 7788 3878
rect 7852 3738 7880 5646
rect 8024 5636 8076 5642
rect 7944 5596 8024 5624
rect 7944 4826 7972 5596
rect 8024 5578 8076 5584
rect 8220 5302 8248 6054
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8404 5302 8432 5578
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8036 4826 8064 4966
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8128 4010 8156 5170
rect 8220 4282 8248 5238
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4282 8340 4558
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8404 4078 8432 5238
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8496 4010 8524 5102
rect 8588 4690 8616 6802
rect 8772 6322 8800 7482
rect 9048 7410 9076 7686
rect 9140 7546 9168 8026
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8864 6322 8892 7346
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8864 6186 8892 6258
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8588 3126 8616 4626
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7760 2582 7788 2858
rect 7852 2650 7880 2994
rect 8680 2854 8708 3470
rect 8956 3398 8984 6938
rect 9048 6322 9076 7346
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6322 9260 6598
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9048 5914 9076 6258
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9232 5778 9260 6258
rect 9324 6236 9352 7822
rect 9416 7478 9444 8434
rect 9692 8430 9720 9472
rect 9876 9432 9904 9998
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10152 9874 10180 10202
rect 10244 9994 10272 10202
rect 10612 10062 10640 11086
rect 11164 10810 11192 11086
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10980 10266 11008 10610
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10060 9738 10088 9862
rect 10152 9846 10272 9874
rect 10060 9710 10180 9738
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9784 9404 9904 9432
rect 9784 8906 9812 9404
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9404 6248 9456 6254
rect 9324 6208 9404 6236
rect 9404 6190 9456 6196
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5166 9444 5510
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4593 9168 4966
rect 9126 4584 9182 4593
rect 9126 4519 9182 4528
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9048 4282 9076 4422
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9140 4146 9168 4519
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9232 4078 9260 4422
rect 9508 4146 9536 8298
rect 9784 7886 9812 8434
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9876 7698 9904 8910
rect 9968 8498 9996 9590
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10060 9178 10088 9522
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9956 8492 10008 8498
rect 10008 8452 10088 8480
rect 9956 8434 10008 8440
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9784 7670 9904 7698
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6798 9720 7142
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 6662 9720 6734
rect 9784 6662 9812 7670
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5914 9628 6054
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9586 5128 9642 5137
rect 9586 5063 9642 5072
rect 9600 5030 9628 5063
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9692 4622 9720 6598
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3126 8984 3334
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 8680 2514 8708 2790
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 9324 2446 9352 3878
rect 9692 3534 9720 3878
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9600 3194 9628 3402
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 32 800 60 2382
rect 940 2372 992 2378
rect 940 2314 992 2320
rect 952 2145 980 2314
rect 938 2136 994 2145
rect 938 2071 994 2080
rect 1964 800 1992 2382
rect 3988 1306 4016 2382
rect 9784 2378 9812 6598
rect 9876 6390 9904 6598
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9968 5234 9996 8298
rect 10060 7886 10088 8452
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10152 7546 10180 9710
rect 10244 9692 10272 9846
rect 10232 9686 10284 9692
rect 10232 9628 10284 9634
rect 10980 9586 11008 10202
rect 11348 10062 11376 11290
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10062 11468 11086
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 10244 9466 10272 9522
rect 10784 9512 10836 9518
rect 10244 9438 10548 9466
rect 10784 9454 10836 9460
rect 10324 9376 10376 9382
rect 10244 9336 10324 9364
rect 10244 9178 10272 9336
rect 10324 9318 10376 9324
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10244 8498 10272 9114
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10336 8673 10364 8774
rect 10322 8664 10378 8673
rect 10322 8599 10378 8608
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10520 8480 10548 9438
rect 10796 9178 10824 9454
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10692 8492 10744 8498
rect 10520 8452 10692 8480
rect 10520 7954 10548 8452
rect 10692 8434 10744 8440
rect 10598 8392 10654 8401
rect 10598 8327 10654 8336
rect 10692 8356 10744 8362
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10612 7750 10640 8327
rect 10692 8298 10744 8304
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10152 6798 10180 7482
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10244 5234 10272 7278
rect 10428 6798 10456 7346
rect 10704 7290 10732 8298
rect 10796 7410 10824 9114
rect 10888 7410 10916 9114
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 8401 11008 8774
rect 11072 8514 11100 9522
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8634 11192 8774
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11072 8486 11192 8514
rect 10966 8392 11022 8401
rect 10966 8327 11022 8336
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10704 7262 10824 7290
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10704 6934 10732 7142
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10336 5166 10364 5782
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10060 4622 10088 5102
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10060 4146 10088 4558
rect 10336 4214 10364 4966
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 9876 3738 9904 4082
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9968 3194 9996 4082
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10060 3126 10088 4082
rect 10152 3738 10180 4082
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10336 3194 10364 3606
rect 10428 3398 10456 6598
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10520 5234 10548 6258
rect 10612 5914 10640 6666
rect 10704 6458 10732 6734
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10796 6322 10824 7262
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10888 6798 10916 6938
rect 10980 6798 11008 8230
rect 11164 7410 11192 8486
rect 11256 8362 11284 9522
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11532 9178 11560 9318
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11520 8968 11572 8974
rect 11334 8936 11390 8945
rect 11520 8910 11572 8916
rect 11334 8871 11390 8880
rect 11348 8362 11376 8871
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10980 6458 11008 6734
rect 11164 6610 11192 7346
rect 11256 6798 11284 7414
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11164 6582 11284 6610
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10612 5234 10640 5578
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10520 4486 10548 5170
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10612 3534 10640 5170
rect 10704 4758 10732 5170
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10796 3942 10824 6258
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5574 11100 6054
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5148 11100 5510
rect 11164 5370 11192 6394
rect 11256 5692 11284 6582
rect 11336 5704 11388 5710
rect 11256 5664 11336 5692
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11256 5302 11284 5664
rect 11336 5646 11388 5652
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11152 5160 11204 5166
rect 11072 5120 11152 5148
rect 11152 5102 11204 5108
rect 11440 4758 11468 7414
rect 11532 7342 11560 8910
rect 11624 8480 11652 10610
rect 11716 9586 11744 11018
rect 11900 9586 11928 15302
rect 13740 12850 13768 15302
rect 14844 15162 14872 15671
rect 15488 15502 15516 17433
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13832 11626 13860 14962
rect 14214 14716 14522 14725
rect 14214 14714 14220 14716
rect 14276 14714 14300 14716
rect 14356 14714 14380 14716
rect 14436 14714 14460 14716
rect 14516 14714 14522 14716
rect 14276 14662 14278 14714
rect 14458 14662 14460 14714
rect 14214 14660 14220 14662
rect 14276 14660 14300 14662
rect 14356 14660 14380 14662
rect 14436 14660 14460 14662
rect 14516 14660 14522 14662
rect 14214 14651 14522 14660
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13924 12170 13952 13874
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14844 13705 14872 13806
rect 14830 13696 14886 13705
rect 14214 13628 14522 13637
rect 14830 13631 14886 13640
rect 14214 13626 14220 13628
rect 14276 13626 14300 13628
rect 14356 13626 14380 13628
rect 14436 13626 14460 13628
rect 14516 13626 14522 13628
rect 14276 13574 14278 13626
rect 14458 13574 14460 13626
rect 14214 13572 14220 13574
rect 14276 13572 14300 13574
rect 14356 13572 14380 13574
rect 14436 13572 14460 13574
rect 14516 13572 14522 13574
rect 14214 13563 14522 13572
rect 14214 12540 14522 12549
rect 14214 12538 14220 12540
rect 14276 12538 14300 12540
rect 14356 12538 14380 12540
rect 14436 12538 14460 12540
rect 14516 12538 14522 12540
rect 14276 12486 14278 12538
rect 14458 12486 14460 12538
rect 14214 12484 14220 12486
rect 14276 12484 14300 12486
rect 14356 12484 14380 12486
rect 14436 12484 14460 12486
rect 14516 12484 14522 12486
rect 14214 12475 14522 12484
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 14214 11452 14522 11461
rect 14214 11450 14220 11452
rect 14276 11450 14300 11452
rect 14356 11450 14380 11452
rect 14436 11450 14460 11452
rect 14516 11450 14522 11452
rect 14276 11398 14278 11450
rect 14458 11398 14460 11450
rect 14214 11396 14220 11398
rect 14276 11396 14300 11398
rect 14356 11396 14380 11398
rect 14436 11396 14460 11398
rect 14516 11396 14522 11398
rect 14214 11387 14522 11396
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14936 10985 14964 11018
rect 14922 10976 14978 10985
rect 14922 10911 14978 10920
rect 14214 10364 14522 10373
rect 14214 10362 14220 10364
rect 14276 10362 14300 10364
rect 14356 10362 14380 10364
rect 14436 10362 14460 10364
rect 14516 10362 14522 10364
rect 14276 10310 14278 10362
rect 14458 10310 14460 10362
rect 14214 10308 14220 10310
rect 14276 10308 14300 10310
rect 14356 10308 14380 10310
rect 14436 10308 14460 10310
rect 14516 10308 14522 10310
rect 14214 10299 14522 10308
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 9042 11928 9522
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11808 8634 11836 8842
rect 11886 8664 11942 8673
rect 11796 8628 11848 8634
rect 11886 8599 11888 8608
rect 11796 8570 11848 8576
rect 11940 8599 11942 8608
rect 11888 8570 11940 8576
rect 11704 8492 11756 8498
rect 11624 8452 11704 8480
rect 11704 8434 11756 8440
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11624 6798 11652 8298
rect 11716 7002 11744 8434
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11532 4826 11560 5578
rect 11624 5030 11652 6734
rect 11808 5710 11836 7686
rect 11992 7410 12020 9930
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12820 8974 12848 9454
rect 14214 9276 14522 9285
rect 14214 9274 14220 9276
rect 14276 9274 14300 9276
rect 14356 9274 14380 9276
rect 14436 9274 14460 9276
rect 14516 9274 14522 9276
rect 14276 9222 14278 9274
rect 14458 9222 14460 9274
rect 14214 9220 14220 9222
rect 14276 9220 14300 9222
rect 14356 9220 14380 9222
rect 14436 9220 14460 9222
rect 14516 9220 14522 9222
rect 14214 9211 14522 9220
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 14462 8936 14518 8945
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8566 12204 8774
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12820 8498 12848 8910
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12820 7954 12848 8434
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 11900 6322 11928 6734
rect 12636 6458 12664 6734
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12820 6322 12848 7890
rect 13280 7750 13308 8910
rect 14462 8871 14518 8880
rect 14476 8566 14504 8871
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14214 8188 14522 8197
rect 14214 8186 14220 8188
rect 14276 8186 14300 8188
rect 14356 8186 14380 8188
rect 14436 8186 14460 8188
rect 14516 8186 14522 8188
rect 14276 8134 14278 8186
rect 14458 8134 14460 8186
rect 14214 8132 14220 8134
rect 14276 8132 14300 8134
rect 14356 8132 14380 8134
rect 14436 8132 14460 8134
rect 14516 8132 14522 8134
rect 14214 8123 14522 8132
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 6798 13308 7686
rect 14214 7100 14522 7109
rect 14214 7098 14220 7100
rect 14276 7098 14300 7100
rect 14356 7098 14380 7100
rect 14436 7098 14460 7100
rect 14516 7098 14522 7100
rect 14276 7046 14278 7098
rect 14458 7046 14460 7098
rect 14214 7044 14220 7046
rect 14276 7044 14300 7046
rect 14356 7044 14380 7046
rect 14436 7044 14460 7046
rect 14516 7044 14522 7046
rect 14214 7035 14522 7044
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12452 5914 12480 6122
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12820 5846 12848 6258
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11428 4752 11480 4758
rect 11480 4700 11560 4706
rect 11428 4694 11560 4700
rect 11440 4678 11560 4694
rect 11532 4622 11560 4678
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11532 4214 11560 4558
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11716 3942 11744 4558
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10520 3058 10548 3402
rect 10612 3058 10640 3470
rect 11716 3466 11744 3878
rect 11808 3738 11836 5646
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12452 5370 12480 5578
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12452 4826 12480 5306
rect 12544 5234 12572 5646
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 12084 3670 12112 4082
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10612 2446 10640 2994
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10796 2514 10824 2790
rect 11072 2650 11100 2994
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11716 2514 11744 3402
rect 12544 3398 12572 5170
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 3058 12572 3334
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 12820 2446 12848 5782
rect 13280 5098 13308 6734
rect 13372 6458 13400 6734
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13372 5370 13400 6394
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14936 6225 14964 6258
rect 14922 6216 14978 6225
rect 14922 6151 14978 6160
rect 14214 6012 14522 6021
rect 14214 6010 14220 6012
rect 14276 6010 14300 6012
rect 14356 6010 14380 6012
rect 14436 6010 14460 6012
rect 14516 6010 14522 6012
rect 14276 5958 14278 6010
rect 14458 5958 14460 6010
rect 14214 5956 14220 5958
rect 14276 5956 14300 5958
rect 14356 5956 14380 5958
rect 14436 5956 14460 5958
rect 14516 5956 14522 5958
rect 14214 5947 14522 5956
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13188 3126 13216 4966
rect 13832 4826 13860 5714
rect 14214 4924 14522 4933
rect 14214 4922 14220 4924
rect 14276 4922 14300 4924
rect 14356 4922 14380 4924
rect 14436 4922 14460 4924
rect 14516 4922 14522 4924
rect 14276 4870 14278 4922
rect 14458 4870 14460 4922
rect 14214 4868 14220 4870
rect 14276 4868 14300 4870
rect 14356 4868 14380 4870
rect 14436 4868 14460 4870
rect 14516 4868 14522 4870
rect 14214 4859 14522 4868
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13924 2446 13952 4218
rect 14936 4185 14964 4422
rect 14922 4176 14978 4185
rect 14922 4111 14978 4120
rect 14214 3836 14522 3845
rect 14214 3834 14220 3836
rect 14276 3834 14300 3836
rect 14356 3834 14380 3836
rect 14436 3834 14460 3836
rect 14516 3834 14522 3836
rect 14276 3782 14278 3834
rect 14458 3782 14460 3834
rect 14214 3780 14220 3782
rect 14276 3780 14300 3782
rect 14356 3780 14380 3782
rect 14436 3780 14460 3782
rect 14516 3780 14522 3782
rect 14214 3771 14522 3780
rect 14214 2748 14522 2757
rect 14214 2746 14220 2748
rect 14276 2746 14300 2748
rect 14356 2746 14380 2748
rect 14436 2746 14460 2748
rect 14516 2746 14522 2748
rect 14276 2694 14278 2746
rect 14458 2694 14460 2746
rect 14214 2692 14220 2694
rect 14276 2692 14300 2694
rect 14356 2692 14380 2694
rect 14436 2692 14460 2694
rect 14516 2692 14522 2694
rect 14214 2683 14522 2692
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 12808 2440 12860 2446
rect 13084 2440 13136 2446
rect 12808 2382 12860 2388
rect 12912 2400 13084 2428
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 3896 1278 4016 1306
rect 3896 800 3924 1278
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 10980 800 11008 2382
rect 12912 800 12940 2400
rect 13084 2382 13136 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14568 1465 14596 2450
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 14554 1456 14610 1465
rect 14554 1391 14610 1400
rect 15488 800 15516 2314
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 15474 0 15530 800
<< via2 >>
rect 938 16360 994 16416
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1398 13640 1454 13696
rect 938 11600 994 11656
rect 938 8900 994 8936
rect 938 8880 940 8900
rect 940 8880 992 8900
rect 992 8880 994 8900
rect 1490 6840 1546 6896
rect 938 4120 994 4176
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 8880 4122 8936
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 5814 9988 5870 10024
rect 5814 9968 5816 9988
rect 5816 9968 5868 9988
rect 5868 9968 5870 9988
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 5722 5072 5778 5128
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5906 3984 5962 4040
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6826 8336 6882 8392
rect 6918 4528 6974 4584
rect 8758 9988 8814 10024
rect 8758 9968 8760 9988
rect 8760 9968 8812 9988
rect 8812 9968 8814 9988
rect 8666 8880 8722 8936
rect 14220 15802 14276 15804
rect 14300 15802 14356 15804
rect 14380 15802 14436 15804
rect 14460 15802 14516 15804
rect 14220 15750 14266 15802
rect 14266 15750 14276 15802
rect 14300 15750 14330 15802
rect 14330 15750 14342 15802
rect 14342 15750 14356 15802
rect 14380 15750 14394 15802
rect 14394 15750 14406 15802
rect 14406 15750 14436 15802
rect 14460 15750 14470 15802
rect 14470 15750 14516 15802
rect 14220 15748 14276 15750
rect 14300 15748 14356 15750
rect 14380 15748 14436 15750
rect 14460 15748 14516 15750
rect 14830 15680 14886 15736
rect 9494 8880 9550 8936
rect 9126 4528 9182 4584
rect 9586 5072 9642 5128
rect 938 2080 994 2136
rect 10322 8608 10378 8664
rect 10598 8336 10654 8392
rect 10966 8336 11022 8392
rect 11334 8880 11390 8936
rect 14220 14714 14276 14716
rect 14300 14714 14356 14716
rect 14380 14714 14436 14716
rect 14460 14714 14516 14716
rect 14220 14662 14266 14714
rect 14266 14662 14276 14714
rect 14300 14662 14330 14714
rect 14330 14662 14342 14714
rect 14342 14662 14356 14714
rect 14380 14662 14394 14714
rect 14394 14662 14406 14714
rect 14406 14662 14436 14714
rect 14460 14662 14470 14714
rect 14470 14662 14516 14714
rect 14220 14660 14276 14662
rect 14300 14660 14356 14662
rect 14380 14660 14436 14662
rect 14460 14660 14516 14662
rect 14830 13640 14886 13696
rect 14220 13626 14276 13628
rect 14300 13626 14356 13628
rect 14380 13626 14436 13628
rect 14460 13626 14516 13628
rect 14220 13574 14266 13626
rect 14266 13574 14276 13626
rect 14300 13574 14330 13626
rect 14330 13574 14342 13626
rect 14342 13574 14356 13626
rect 14380 13574 14394 13626
rect 14394 13574 14406 13626
rect 14406 13574 14436 13626
rect 14460 13574 14470 13626
rect 14470 13574 14516 13626
rect 14220 13572 14276 13574
rect 14300 13572 14356 13574
rect 14380 13572 14436 13574
rect 14460 13572 14516 13574
rect 14220 12538 14276 12540
rect 14300 12538 14356 12540
rect 14380 12538 14436 12540
rect 14460 12538 14516 12540
rect 14220 12486 14266 12538
rect 14266 12486 14276 12538
rect 14300 12486 14330 12538
rect 14330 12486 14342 12538
rect 14342 12486 14356 12538
rect 14380 12486 14394 12538
rect 14394 12486 14406 12538
rect 14406 12486 14436 12538
rect 14460 12486 14470 12538
rect 14470 12486 14516 12538
rect 14220 12484 14276 12486
rect 14300 12484 14356 12486
rect 14380 12484 14436 12486
rect 14460 12484 14516 12486
rect 14220 11450 14276 11452
rect 14300 11450 14356 11452
rect 14380 11450 14436 11452
rect 14460 11450 14516 11452
rect 14220 11398 14266 11450
rect 14266 11398 14276 11450
rect 14300 11398 14330 11450
rect 14330 11398 14342 11450
rect 14342 11398 14356 11450
rect 14380 11398 14394 11450
rect 14394 11398 14406 11450
rect 14406 11398 14436 11450
rect 14460 11398 14470 11450
rect 14470 11398 14516 11450
rect 14220 11396 14276 11398
rect 14300 11396 14356 11398
rect 14380 11396 14436 11398
rect 14460 11396 14516 11398
rect 14922 10920 14978 10976
rect 14220 10362 14276 10364
rect 14300 10362 14356 10364
rect 14380 10362 14436 10364
rect 14460 10362 14516 10364
rect 14220 10310 14266 10362
rect 14266 10310 14276 10362
rect 14300 10310 14330 10362
rect 14330 10310 14342 10362
rect 14342 10310 14356 10362
rect 14380 10310 14394 10362
rect 14394 10310 14406 10362
rect 14406 10310 14436 10362
rect 14460 10310 14470 10362
rect 14470 10310 14516 10362
rect 14220 10308 14276 10310
rect 14300 10308 14356 10310
rect 14380 10308 14436 10310
rect 14460 10308 14516 10310
rect 11886 8628 11942 8664
rect 11886 8608 11888 8628
rect 11888 8608 11940 8628
rect 11940 8608 11942 8628
rect 14220 9274 14276 9276
rect 14300 9274 14356 9276
rect 14380 9274 14436 9276
rect 14460 9274 14516 9276
rect 14220 9222 14266 9274
rect 14266 9222 14276 9274
rect 14300 9222 14330 9274
rect 14330 9222 14342 9274
rect 14342 9222 14356 9274
rect 14380 9222 14394 9274
rect 14394 9222 14406 9274
rect 14406 9222 14436 9274
rect 14460 9222 14470 9274
rect 14470 9222 14516 9274
rect 14220 9220 14276 9222
rect 14300 9220 14356 9222
rect 14380 9220 14436 9222
rect 14460 9220 14516 9222
rect 14462 8880 14518 8936
rect 14220 8186 14276 8188
rect 14300 8186 14356 8188
rect 14380 8186 14436 8188
rect 14460 8186 14516 8188
rect 14220 8134 14266 8186
rect 14266 8134 14276 8186
rect 14300 8134 14330 8186
rect 14330 8134 14342 8186
rect 14342 8134 14356 8186
rect 14380 8134 14394 8186
rect 14394 8134 14406 8186
rect 14406 8134 14436 8186
rect 14460 8134 14470 8186
rect 14470 8134 14516 8186
rect 14220 8132 14276 8134
rect 14300 8132 14356 8134
rect 14380 8132 14436 8134
rect 14460 8132 14516 8134
rect 14220 7098 14276 7100
rect 14300 7098 14356 7100
rect 14380 7098 14436 7100
rect 14460 7098 14516 7100
rect 14220 7046 14266 7098
rect 14266 7046 14276 7098
rect 14300 7046 14330 7098
rect 14330 7046 14342 7098
rect 14342 7046 14356 7098
rect 14380 7046 14394 7098
rect 14394 7046 14406 7098
rect 14406 7046 14436 7098
rect 14460 7046 14470 7098
rect 14470 7046 14516 7098
rect 14220 7044 14276 7046
rect 14300 7044 14356 7046
rect 14380 7044 14436 7046
rect 14460 7044 14516 7046
rect 14922 6160 14978 6216
rect 14220 6010 14276 6012
rect 14300 6010 14356 6012
rect 14380 6010 14436 6012
rect 14460 6010 14516 6012
rect 14220 5958 14266 6010
rect 14266 5958 14276 6010
rect 14300 5958 14330 6010
rect 14330 5958 14342 6010
rect 14342 5958 14356 6010
rect 14380 5958 14394 6010
rect 14394 5958 14406 6010
rect 14406 5958 14436 6010
rect 14460 5958 14470 6010
rect 14470 5958 14516 6010
rect 14220 5956 14276 5958
rect 14300 5956 14356 5958
rect 14380 5956 14436 5958
rect 14460 5956 14516 5958
rect 14220 4922 14276 4924
rect 14300 4922 14356 4924
rect 14380 4922 14436 4924
rect 14460 4922 14516 4924
rect 14220 4870 14266 4922
rect 14266 4870 14276 4922
rect 14300 4870 14330 4922
rect 14330 4870 14342 4922
rect 14342 4870 14356 4922
rect 14380 4870 14394 4922
rect 14394 4870 14406 4922
rect 14406 4870 14436 4922
rect 14460 4870 14470 4922
rect 14470 4870 14516 4922
rect 14220 4868 14276 4870
rect 14300 4868 14356 4870
rect 14380 4868 14436 4870
rect 14460 4868 14516 4870
rect 14922 4120 14978 4176
rect 14220 3834 14276 3836
rect 14300 3834 14356 3836
rect 14380 3834 14436 3836
rect 14460 3834 14516 3836
rect 14220 3782 14266 3834
rect 14266 3782 14276 3834
rect 14300 3782 14330 3834
rect 14330 3782 14342 3834
rect 14342 3782 14356 3834
rect 14380 3782 14394 3834
rect 14394 3782 14406 3834
rect 14406 3782 14436 3834
rect 14460 3782 14470 3834
rect 14470 3782 14516 3834
rect 14220 3780 14276 3782
rect 14300 3780 14356 3782
rect 14380 3780 14436 3782
rect 14460 3780 14516 3782
rect 14220 2746 14276 2748
rect 14300 2746 14356 2748
rect 14380 2746 14436 2748
rect 14460 2746 14516 2748
rect 14220 2694 14266 2746
rect 14266 2694 14276 2746
rect 14300 2694 14330 2746
rect 14330 2694 14342 2746
rect 14342 2694 14356 2746
rect 14380 2694 14394 2746
rect 14394 2694 14406 2746
rect 14406 2694 14436 2746
rect 14460 2694 14470 2746
rect 14470 2694 14516 2746
rect 14220 2692 14276 2694
rect 14300 2692 14356 2694
rect 14380 2692 14436 2694
rect 14460 2692 14516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 14554 1400 14610 1456
<< metal3 >>
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 14210 15808 14526 15809
rect 14210 15744 14216 15808
rect 14280 15744 14296 15808
rect 14360 15744 14376 15808
rect 14440 15744 14456 15808
rect 14520 15744 14526 15808
rect 14210 15743 14526 15744
rect 14825 15738 14891 15741
rect 15289 15738 16089 15768
rect 14825 15736 16089 15738
rect 14825 15680 14830 15736
rect 14886 15680 16089 15736
rect 14825 15678 16089 15680
rect 14825 15675 14891 15678
rect 15289 15648 16089 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 14210 14720 14526 14721
rect 14210 14656 14216 14720
rect 14280 14656 14296 14720
rect 14360 14656 14376 14720
rect 14440 14656 14456 14720
rect 14520 14656 14526 14720
rect 14210 14655 14526 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 14825 13698 14891 13701
rect 15289 13698 16089 13728
rect 14825 13696 16089 13698
rect 14825 13640 14830 13696
rect 14886 13640 16089 13696
rect 14825 13638 16089 13640
rect 14825 13635 14891 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 14210 13632 14526 13633
rect 14210 13568 14216 13632
rect 14280 13568 14296 13632
rect 14360 13568 14376 13632
rect 14440 13568 14456 13632
rect 14520 13568 14526 13632
rect 15289 13608 16089 13638
rect 14210 13567 14526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 14210 12544 14526 12545
rect 14210 12480 14216 12544
rect 14280 12480 14296 12544
rect 14360 12480 14376 12544
rect 14440 12480 14456 12544
rect 14520 12480 14526 12544
rect 14210 12479 14526 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 14210 11456 14526 11457
rect 14210 11392 14216 11456
rect 14280 11392 14296 11456
rect 14360 11392 14376 11456
rect 14440 11392 14456 11456
rect 14520 11392 14526 11456
rect 14210 11391 14526 11392
rect 14917 10978 14983 10981
rect 15289 10978 16089 11008
rect 14917 10976 16089 10978
rect 14917 10920 14922 10976
rect 14978 10920 16089 10976
rect 14917 10918 16089 10920
rect 14917 10915 14983 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 15289 10888 16089 10918
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 14210 10368 14526 10369
rect 14210 10304 14216 10368
rect 14280 10304 14296 10368
rect 14360 10304 14376 10368
rect 14440 10304 14456 10368
rect 14520 10304 14526 10368
rect 14210 10303 14526 10304
rect 5809 10026 5875 10029
rect 8753 10026 8819 10029
rect 5809 10024 8819 10026
rect 5809 9968 5814 10024
rect 5870 9968 8758 10024
rect 8814 9968 8819 10024
rect 5809 9966 8819 9968
rect 5809 9963 5875 9966
rect 8753 9963 8819 9966
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 14210 9280 14526 9281
rect 14210 9216 14216 9280
rect 14280 9216 14296 9280
rect 14360 9216 14376 9280
rect 14440 9216 14456 9280
rect 14520 9216 14526 9280
rect 14210 9215 14526 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 4061 8938 4127 8941
rect 8661 8938 8727 8941
rect 4061 8936 8727 8938
rect 4061 8880 4066 8936
rect 4122 8880 8666 8936
rect 8722 8880 8727 8936
rect 4061 8878 8727 8880
rect 4061 8875 4127 8878
rect 8661 8875 8727 8878
rect 9489 8938 9555 8941
rect 11329 8938 11395 8941
rect 9489 8936 11395 8938
rect 9489 8880 9494 8936
rect 9550 8880 11334 8936
rect 11390 8880 11395 8936
rect 9489 8878 11395 8880
rect 9489 8875 9555 8878
rect 11329 8875 11395 8878
rect 14457 8938 14523 8941
rect 15289 8938 16089 8968
rect 14457 8936 16089 8938
rect 14457 8880 14462 8936
rect 14518 8880 16089 8936
rect 14457 8878 16089 8880
rect 14457 8875 14523 8878
rect 15289 8848 16089 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 10317 8666 10383 8669
rect 11881 8666 11947 8669
rect 10317 8664 11947 8666
rect 10317 8608 10322 8664
rect 10378 8608 11886 8664
rect 11942 8608 11947 8664
rect 10317 8606 11947 8608
rect 10317 8603 10383 8606
rect 11881 8603 11947 8606
rect 6821 8396 6887 8397
rect 6821 8394 6868 8396
rect 6776 8392 6868 8394
rect 6776 8336 6826 8392
rect 6776 8334 6868 8336
rect 6821 8332 6868 8334
rect 6932 8332 6938 8396
rect 10593 8394 10659 8397
rect 10961 8394 11027 8397
rect 10593 8392 11027 8394
rect 10593 8336 10598 8392
rect 10654 8336 10966 8392
rect 11022 8336 11027 8392
rect 10593 8334 11027 8336
rect 6821 8331 6887 8332
rect 10593 8331 10659 8334
rect 10961 8331 11027 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 14210 8192 14526 8193
rect 14210 8128 14216 8192
rect 14280 8128 14296 8192
rect 14360 8128 14376 8192
rect 14440 8128 14456 8192
rect 14520 8128 14526 8192
rect 14210 8127 14526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 14210 7104 14526 7105
rect 14210 7040 14216 7104
rect 14280 7040 14296 7104
rect 14360 7040 14376 7104
rect 14440 7040 14456 7104
rect 14520 7040 14526 7104
rect 14210 7039 14526 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 14917 6218 14983 6221
rect 15289 6218 16089 6248
rect 14917 6216 16089 6218
rect 14917 6160 14922 6216
rect 14978 6160 16089 6216
rect 14917 6158 16089 6160
rect 14917 6155 14983 6158
rect 15289 6128 16089 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 14210 6016 14526 6017
rect 14210 5952 14216 6016
rect 14280 5952 14296 6016
rect 14360 5952 14376 6016
rect 14440 5952 14456 6016
rect 14520 5952 14526 6016
rect 14210 5951 14526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 5717 5130 5783 5133
rect 9581 5130 9647 5133
rect 5717 5128 9647 5130
rect 5717 5072 5722 5128
rect 5778 5072 9586 5128
rect 9642 5072 9647 5128
rect 5717 5070 9647 5072
rect 5717 5067 5783 5070
rect 9581 5067 9647 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 14210 4928 14526 4929
rect 14210 4864 14216 4928
rect 14280 4864 14296 4928
rect 14360 4864 14376 4928
rect 14440 4864 14456 4928
rect 14520 4864 14526 4928
rect 14210 4863 14526 4864
rect 6913 4586 6979 4589
rect 9121 4586 9187 4589
rect 6913 4584 9187 4586
rect 6913 4528 6918 4584
rect 6974 4528 9126 4584
rect 9182 4528 9187 4584
rect 6913 4526 9187 4528
rect 6913 4523 6979 4526
rect 9121 4523 9187 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 14917 4178 14983 4181
rect 15289 4178 16089 4208
rect 14917 4176 16089 4178
rect 14917 4120 14922 4176
rect 14978 4120 16089 4176
rect 14917 4118 16089 4120
rect 14917 4115 14983 4118
rect 15289 4088 16089 4118
rect 5901 4042 5967 4045
rect 6862 4042 6868 4044
rect 5901 4040 6868 4042
rect 5901 3984 5906 4040
rect 5962 3984 6868 4040
rect 5901 3982 6868 3984
rect 5901 3979 5967 3982
rect 6862 3980 6868 3982
rect 6932 3980 6938 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 14210 3840 14526 3841
rect 14210 3776 14216 3840
rect 14280 3776 14296 3840
rect 14360 3776 14376 3840
rect 14440 3776 14456 3840
rect 14520 3776 14526 3840
rect 14210 3775 14526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 14210 2752 14526 2753
rect 14210 2688 14216 2752
rect 14280 2688 14296 2752
rect 14360 2688 14376 2752
rect 14440 2688 14456 2752
rect 14520 2688 14526 2752
rect 14210 2687 14526 2688
rect 4870 2208 5186 2209
rect 0 2138 800 2168
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 933 2138 999 2141
rect 0 2136 999 2138
rect 0 2080 938 2136
rect 994 2080 999 2136
rect 0 2078 999 2080
rect 0 2048 800 2078
rect 933 2075 999 2078
rect 14549 1458 14615 1461
rect 15289 1458 16089 1488
rect 14549 1456 16089 1458
rect 14549 1400 14554 1456
rect 14610 1400 16089 1456
rect 14549 1398 16089 1400
rect 14549 1395 14615 1398
rect 15289 1368 16089 1398
<< via3 >>
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 14216 15804 14280 15808
rect 14216 15748 14220 15804
rect 14220 15748 14276 15804
rect 14276 15748 14280 15804
rect 14216 15744 14280 15748
rect 14296 15804 14360 15808
rect 14296 15748 14300 15804
rect 14300 15748 14356 15804
rect 14356 15748 14360 15804
rect 14296 15744 14360 15748
rect 14376 15804 14440 15808
rect 14376 15748 14380 15804
rect 14380 15748 14436 15804
rect 14436 15748 14440 15804
rect 14376 15744 14440 15748
rect 14456 15804 14520 15808
rect 14456 15748 14460 15804
rect 14460 15748 14516 15804
rect 14516 15748 14520 15804
rect 14456 15744 14520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 14216 14716 14280 14720
rect 14216 14660 14220 14716
rect 14220 14660 14276 14716
rect 14276 14660 14280 14716
rect 14216 14656 14280 14660
rect 14296 14716 14360 14720
rect 14296 14660 14300 14716
rect 14300 14660 14356 14716
rect 14356 14660 14360 14716
rect 14296 14656 14360 14660
rect 14376 14716 14440 14720
rect 14376 14660 14380 14716
rect 14380 14660 14436 14716
rect 14436 14660 14440 14716
rect 14376 14656 14440 14660
rect 14456 14716 14520 14720
rect 14456 14660 14460 14716
rect 14460 14660 14516 14716
rect 14516 14660 14520 14716
rect 14456 14656 14520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 14216 13628 14280 13632
rect 14216 13572 14220 13628
rect 14220 13572 14276 13628
rect 14276 13572 14280 13628
rect 14216 13568 14280 13572
rect 14296 13628 14360 13632
rect 14296 13572 14300 13628
rect 14300 13572 14356 13628
rect 14356 13572 14360 13628
rect 14296 13568 14360 13572
rect 14376 13628 14440 13632
rect 14376 13572 14380 13628
rect 14380 13572 14436 13628
rect 14436 13572 14440 13628
rect 14376 13568 14440 13572
rect 14456 13628 14520 13632
rect 14456 13572 14460 13628
rect 14460 13572 14516 13628
rect 14516 13572 14520 13628
rect 14456 13568 14520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 14216 12540 14280 12544
rect 14216 12484 14220 12540
rect 14220 12484 14276 12540
rect 14276 12484 14280 12540
rect 14216 12480 14280 12484
rect 14296 12540 14360 12544
rect 14296 12484 14300 12540
rect 14300 12484 14356 12540
rect 14356 12484 14360 12540
rect 14296 12480 14360 12484
rect 14376 12540 14440 12544
rect 14376 12484 14380 12540
rect 14380 12484 14436 12540
rect 14436 12484 14440 12540
rect 14376 12480 14440 12484
rect 14456 12540 14520 12544
rect 14456 12484 14460 12540
rect 14460 12484 14516 12540
rect 14516 12484 14520 12540
rect 14456 12480 14520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 14216 11452 14280 11456
rect 14216 11396 14220 11452
rect 14220 11396 14276 11452
rect 14276 11396 14280 11452
rect 14216 11392 14280 11396
rect 14296 11452 14360 11456
rect 14296 11396 14300 11452
rect 14300 11396 14356 11452
rect 14356 11396 14360 11452
rect 14296 11392 14360 11396
rect 14376 11452 14440 11456
rect 14376 11396 14380 11452
rect 14380 11396 14436 11452
rect 14436 11396 14440 11452
rect 14376 11392 14440 11396
rect 14456 11452 14520 11456
rect 14456 11396 14460 11452
rect 14460 11396 14516 11452
rect 14516 11396 14520 11452
rect 14456 11392 14520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 14216 10364 14280 10368
rect 14216 10308 14220 10364
rect 14220 10308 14276 10364
rect 14276 10308 14280 10364
rect 14216 10304 14280 10308
rect 14296 10364 14360 10368
rect 14296 10308 14300 10364
rect 14300 10308 14356 10364
rect 14356 10308 14360 10364
rect 14296 10304 14360 10308
rect 14376 10364 14440 10368
rect 14376 10308 14380 10364
rect 14380 10308 14436 10364
rect 14436 10308 14440 10364
rect 14376 10304 14440 10308
rect 14456 10364 14520 10368
rect 14456 10308 14460 10364
rect 14460 10308 14516 10364
rect 14516 10308 14520 10364
rect 14456 10304 14520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 14216 9276 14280 9280
rect 14216 9220 14220 9276
rect 14220 9220 14276 9276
rect 14276 9220 14280 9276
rect 14216 9216 14280 9220
rect 14296 9276 14360 9280
rect 14296 9220 14300 9276
rect 14300 9220 14356 9276
rect 14356 9220 14360 9276
rect 14296 9216 14360 9220
rect 14376 9276 14440 9280
rect 14376 9220 14380 9276
rect 14380 9220 14436 9276
rect 14436 9220 14440 9276
rect 14376 9216 14440 9220
rect 14456 9276 14520 9280
rect 14456 9220 14460 9276
rect 14460 9220 14516 9276
rect 14516 9220 14520 9276
rect 14456 9216 14520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 6868 8392 6932 8396
rect 6868 8336 6882 8392
rect 6882 8336 6932 8392
rect 6868 8332 6932 8336
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 14216 8188 14280 8192
rect 14216 8132 14220 8188
rect 14220 8132 14276 8188
rect 14276 8132 14280 8188
rect 14216 8128 14280 8132
rect 14296 8188 14360 8192
rect 14296 8132 14300 8188
rect 14300 8132 14356 8188
rect 14356 8132 14360 8188
rect 14296 8128 14360 8132
rect 14376 8188 14440 8192
rect 14376 8132 14380 8188
rect 14380 8132 14436 8188
rect 14436 8132 14440 8188
rect 14376 8128 14440 8132
rect 14456 8188 14520 8192
rect 14456 8132 14460 8188
rect 14460 8132 14516 8188
rect 14516 8132 14520 8188
rect 14456 8128 14520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 14216 7100 14280 7104
rect 14216 7044 14220 7100
rect 14220 7044 14276 7100
rect 14276 7044 14280 7100
rect 14216 7040 14280 7044
rect 14296 7100 14360 7104
rect 14296 7044 14300 7100
rect 14300 7044 14356 7100
rect 14356 7044 14360 7100
rect 14296 7040 14360 7044
rect 14376 7100 14440 7104
rect 14376 7044 14380 7100
rect 14380 7044 14436 7100
rect 14436 7044 14440 7100
rect 14376 7040 14440 7044
rect 14456 7100 14520 7104
rect 14456 7044 14460 7100
rect 14460 7044 14516 7100
rect 14516 7044 14520 7100
rect 14456 7040 14520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 14216 6012 14280 6016
rect 14216 5956 14220 6012
rect 14220 5956 14276 6012
rect 14276 5956 14280 6012
rect 14216 5952 14280 5956
rect 14296 6012 14360 6016
rect 14296 5956 14300 6012
rect 14300 5956 14356 6012
rect 14356 5956 14360 6012
rect 14296 5952 14360 5956
rect 14376 6012 14440 6016
rect 14376 5956 14380 6012
rect 14380 5956 14436 6012
rect 14436 5956 14440 6012
rect 14376 5952 14440 5956
rect 14456 6012 14520 6016
rect 14456 5956 14460 6012
rect 14460 5956 14516 6012
rect 14516 5956 14520 6012
rect 14456 5952 14520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 14216 4924 14280 4928
rect 14216 4868 14220 4924
rect 14220 4868 14276 4924
rect 14276 4868 14280 4924
rect 14216 4864 14280 4868
rect 14296 4924 14360 4928
rect 14296 4868 14300 4924
rect 14300 4868 14356 4924
rect 14356 4868 14360 4924
rect 14296 4864 14360 4868
rect 14376 4924 14440 4928
rect 14376 4868 14380 4924
rect 14380 4868 14436 4924
rect 14436 4868 14440 4924
rect 14376 4864 14440 4868
rect 14456 4924 14520 4928
rect 14456 4868 14460 4924
rect 14460 4868 14516 4924
rect 14516 4868 14520 4924
rect 14456 4864 14520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 6868 3980 6932 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 14216 3836 14280 3840
rect 14216 3780 14220 3836
rect 14220 3780 14276 3836
rect 14276 3780 14280 3836
rect 14216 3776 14280 3780
rect 14296 3836 14360 3840
rect 14296 3780 14300 3836
rect 14300 3780 14356 3836
rect 14356 3780 14360 3836
rect 14296 3776 14360 3780
rect 14376 3836 14440 3840
rect 14376 3780 14380 3836
rect 14380 3780 14436 3836
rect 14436 3780 14440 3836
rect 14376 3776 14440 3780
rect 14456 3836 14520 3840
rect 14456 3780 14460 3836
rect 14460 3780 14516 3836
rect 14516 3780 14520 3836
rect 14456 3776 14520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 14216 2748 14280 2752
rect 14216 2692 14220 2748
rect 14220 2692 14276 2748
rect 14276 2692 14280 2748
rect 14216 2688 14280 2692
rect 14296 2748 14360 2752
rect 14296 2692 14300 2748
rect 14300 2692 14356 2748
rect 14356 2692 14360 2748
rect 14296 2688 14360 2692
rect 14376 2748 14440 2752
rect 14376 2692 14380 2748
rect 14380 2692 14436 2748
rect 14436 2692 14440 2748
rect 14376 2688 14440 2692
rect 14456 2748 14520 2752
rect 14456 2692 14460 2748
rect 14460 2692 14516 2748
rect 14516 2692 14520 2748
rect 14456 2688 14520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 15808 4528 15824
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15624 4528 15744
rect 4208 15388 4250 15624
rect 4486 15388 4528 15624
rect 4208 14720 4528 15388
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 15264 5188 15824
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 14208 15808 14528 15824
rect 14208 15744 14216 15808
rect 14280 15744 14296 15808
rect 14360 15744 14376 15808
rect 14440 15744 14456 15808
rect 14520 15744 14528 15808
rect 14208 15624 14528 15744
rect 14208 15388 14250 15624
rect 14486 15388 14528 15624
rect 14208 14720 14528 15388
rect 14208 14656 14216 14720
rect 14280 14656 14296 14720
rect 14360 14656 14376 14720
rect 14440 14656 14456 14720
rect 14520 14656 14528 14720
rect 14208 13632 14528 14656
rect 14208 13568 14216 13632
rect 14280 13568 14296 13632
rect 14360 13568 14376 13632
rect 14440 13568 14456 13632
rect 14520 13568 14528 13632
rect 14208 12544 14528 13568
rect 14208 12480 14216 12544
rect 14280 12480 14296 12544
rect 14360 12480 14376 12544
rect 14440 12480 14456 12544
rect 14520 12480 14528 12544
rect 14208 11456 14528 12480
rect 14208 11392 14216 11456
rect 14280 11392 14296 11456
rect 14360 11392 14376 11456
rect 14440 11392 14456 11456
rect 14520 11392 14528 11456
rect 14208 10368 14528 11392
rect 14208 10304 14216 10368
rect 14280 10304 14296 10368
rect 14360 10304 14376 10368
rect 14440 10304 14456 10368
rect 14520 10304 14528 10368
rect 14208 9280 14528 10304
rect 14208 9216 14216 9280
rect 14280 9216 14296 9280
rect 14360 9216 14376 9280
rect 14440 9216 14456 9280
rect 14520 9216 14528 9280
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 6870 4045 6930 8331
rect 14208 8192 14528 9216
rect 14208 8128 14216 8192
rect 14280 8128 14296 8192
rect 14360 8128 14376 8192
rect 14440 8128 14456 8192
rect 14520 8128 14528 8192
rect 14208 7104 14528 8128
rect 14208 7040 14216 7104
rect 14280 7040 14296 7104
rect 14360 7040 14376 7104
rect 14440 7040 14456 7104
rect 14520 7040 14528 7104
rect 14208 6016 14528 7040
rect 14208 5952 14216 6016
rect 14280 5952 14296 6016
rect 14360 5952 14376 6016
rect 14440 5952 14456 6016
rect 14520 5952 14528 6016
rect 14208 5624 14528 5952
rect 14208 5388 14250 5624
rect 14486 5388 14528 5624
rect 14208 4928 14528 5388
rect 14208 4864 14216 4928
rect 14280 4864 14296 4928
rect 14360 4864 14376 4928
rect 14440 4864 14456 4928
rect 14520 4864 14528 4928
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 14208 3840 14528 4864
rect 14208 3776 14216 3840
rect 14280 3776 14296 3840
rect 14360 3776 14376 3840
rect 14440 3776 14456 3840
rect 14520 3776 14528 3840
rect 14208 2752 14528 3776
rect 14208 2688 14216 2752
rect 14280 2688 14296 2752
rect 14360 2688 14376 2752
rect 14440 2688 14456 2752
rect 14520 2688 14528 2752
rect 14208 2128 14528 2688
<< via4 >>
rect 4250 15388 4486 15624
rect 4250 5388 4486 5624
rect 14250 15388 14486 15624
rect 14250 5388 14486 5624
<< metal5 >>
rect 1056 15624 14952 15666
rect 1056 15388 4250 15624
rect 4486 15388 14250 15624
rect 14486 15388 14952 15624
rect 1056 15346 14952 15388
rect 1056 5624 14952 5666
rect 1056 5388 4250 5624
rect 4486 5388 14250 5624
rect 14486 5388 14952 5624
rect 1056 5346 14952 5388
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 0
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _151_
timestamp 0
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _152_
timestamp 0
transform -1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _153_
timestamp 0
transform 1 0 4600 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 0
transform -1 0 3128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 0
transform -1 0 3680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _156_
timestamp 0
transform 1 0 3956 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _157_
timestamp 0
transform -1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _158_
timestamp 0
transform -1 0 5888 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _159_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _160_
timestamp 0
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _161_
timestamp 0
transform 1 0 3496 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_4  _162_
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _163_
timestamp 0
transform -1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _164_
timestamp 0
transform 1 0 4416 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _165_
timestamp 0
transform 1 0 11684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _166_
timestamp 0
transform -1 0 12788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _167_
timestamp 0
transform -1 0 12788 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _168_
timestamp 0
transform -1 0 13432 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _169_
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _170_
timestamp 0
transform 1 0 4968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _171_
timestamp 0
transform 1 0 6716 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _172_
timestamp 0
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _173_
timestamp 0
transform -1 0 10580 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _174_
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _175_
timestamp 0
transform -1 0 8464 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _176_
timestamp 0
transform -1 0 13524 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _177_
timestamp 0
transform 1 0 6072 0 1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _178_
timestamp 0
transform 1 0 3496 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _179_
timestamp 0
transform 1 0 4232 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _180_
timestamp 0
transform -1 0 5244 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _181_
timestamp 0
transform -1 0 4876 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 0
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _183_
timestamp 0
transform -1 0 10948 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _184_
timestamp 0
transform 1 0 9660 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _185_
timestamp 0
transform 1 0 8096 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _186_
timestamp 0
transform 1 0 9292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 0
transform -1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 0
transform 1 0 12788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _189_
timestamp 0
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _190_
timestamp 0
transform -1 0 12144 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _191_
timestamp 0
transform -1 0 9384 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _192_
timestamp 0
transform -1 0 8280 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _193_
timestamp 0
transform 1 0 5060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _194_
timestamp 0
transform 1 0 4784 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _195_
timestamp 0
transform -1 0 5336 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _196_
timestamp 0
transform 1 0 7544 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _197_
timestamp 0
transform -1 0 8648 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _198_
timestamp 0
transform -1 0 7084 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _199_
timestamp 0
transform 1 0 5336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _200_
timestamp 0
transform 1 0 6072 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2o_4  _201_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__or3_4  _202_
timestamp 0
transform -1 0 7176 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _203_
timestamp 0
transform 1 0 6532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _204_
timestamp 0
transform 1 0 4600 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _205_
timestamp 0
transform 1 0 5336 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _206_
timestamp 0
transform -1 0 7636 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 0
transform 1 0 5336 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _208_
timestamp 0
transform 1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _209_
timestamp 0
transform 1 0 6072 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _210_
timestamp 0
transform 1 0 3956 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _211_
timestamp 0
transform -1 0 4232 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2o_1  _212_
timestamp 0
transform 1 0 3680 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _213_
timestamp 0
transform 1 0 4048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _214_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _215_
timestamp 0
transform 1 0 2760 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _216_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 0
transform -1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _218_
timestamp 0
transform -1 0 5152 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _219_
timestamp 0
transform -1 0 6256 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _220_
timestamp 0
transform -1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _221_
timestamp 0
transform -1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _222_
timestamp 0
transform 1 0 7084 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _223_
timestamp 0
transform 1 0 6348 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _224_
timestamp 0
transform 1 0 5612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _225_
timestamp 0
transform 1 0 6440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _226_
timestamp 0
transform 1 0 6992 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _227_
timestamp 0
transform 1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _228_
timestamp 0
transform 1 0 7820 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _229_
timestamp 0
transform 1 0 6440 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _230_
timestamp 0
transform -1 0 7820 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _231_
timestamp 0
transform -1 0 8648 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _232_
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _233_
timestamp 0
transform -1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _234_
timestamp 0
transform -1 0 11500 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 0
transform -1 0 11316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _236_
timestamp 0
transform 1 0 10856 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _237_
timestamp 0
transform 1 0 10304 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _238_
timestamp 0
transform -1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _239_
timestamp 0
transform 1 0 9016 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _240_
timestamp 0
transform 1 0 9108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _241_
timestamp 0
transform 1 0 8924 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _242_
timestamp 0
transform 1 0 9200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _243_
timestamp 0
transform 1 0 9200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _244_
timestamp 0
transform 1 0 9568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _245_
timestamp 0
transform 1 0 10580 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _246_
timestamp 0
transform -1 0 11316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _247_
timestamp 0
transform -1 0 13340 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__o211a_1  _248_
timestamp 0
transform 1 0 10120 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 0
transform 1 0 10304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _250_
timestamp 0
transform -1 0 8464 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _251_
timestamp 0
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _252_
timestamp 0
transform 1 0 9384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _253_
timestamp 0
transform 1 0 7912 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _254_
timestamp 0
transform -1 0 9200 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _255_
timestamp 0
transform 1 0 8096 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _256_
timestamp 0
transform 1 0 10672 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _257_
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _258_
timestamp 0
transform -1 0 12144 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _259_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _260_
timestamp 0
transform -1 0 11868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _261_
timestamp 0
transform 1 0 8924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _262_
timestamp 0
transform 1 0 9476 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _263_
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _265_
timestamp 0
transform 1 0 12880 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _266_
timestamp 0
transform -1 0 12880 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _267_
timestamp 0
transform -1 0 11684 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _268_
timestamp 0
transform -1 0 11776 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _269_
timestamp 0
transform -1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _270_
timestamp 0
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _271_
timestamp 0
transform -1 0 12144 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _272_
timestamp 0
transform 1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _273_
timestamp 0
transform 1 0 10672 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _274_
timestamp 0
transform -1 0 12236 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _275_
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _276_
timestamp 0
transform -1 0 12052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _277_
timestamp 0
transform -1 0 13156 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _278_
timestamp 0
transform 1 0 8648 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _279_
timestamp 0
transform 1 0 7912 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _280_
timestamp 0
transform 1 0 7912 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _281_
timestamp 0
transform 1 0 9384 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _282_
timestamp 0
transform -1 0 10580 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _283_
timestamp 0
transform 1 0 9936 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _284_
timestamp 0
transform -1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _285_
timestamp 0
transform 1 0 8924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _286_
timestamp 0
transform 1 0 9568 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _287_
timestamp 0
transform 1 0 10212 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _288_
timestamp 0
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _289_
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _290_
timestamp 0
transform 1 0 8924 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _291_
timestamp 0
transform 1 0 7820 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _292_
timestamp 0
transform -1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _293_
timestamp 0
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _294_
timestamp 0
transform 1 0 6440 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _295_
timestamp 0
transform -1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _296_
timestamp 0
transform -1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _297_
timestamp 0
transform -1 0 8832 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _298_
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _299_
timestamp 0
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _300_
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _301_
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _303_
timestamp 0
transform 1 0 5520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _304_
timestamp 0
transform -1 0 6164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _305_
timestamp 0
transform -1 0 8004 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _306_
timestamp 0
transform 1 0 7544 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _307_
timestamp 0
transform -1 0 10488 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__a31oi_1  _308_
timestamp 0
transform 1 0 6256 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _309_
timestamp 0
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_16
timestamp 0
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 0
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_63
timestamp 0
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_77
timestamp 0
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_90
timestamp 0
transform 1 0 9384 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_102
timestamp 0
transform 1 0 10488 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 0
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_65
timestamp 0
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_84
timestamp 0
transform 1 0 8832 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_91
timestamp 0
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 0
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_120
timestamp 0
transform 1 0 12144 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_132
timestamp 0
transform 1 0 13248 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_144
timestamp 0
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_59
timestamp 0
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_71
timestamp 0
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_78
timestamp 0
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 0
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_107
timestamp 0
transform 1 0 10948 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_50
timestamp 0
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_73
timestamp 0
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_92
timestamp 0
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_100
timestamp 0
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_119
timestamp 0
transform 1 0 12052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_131
timestamp 0
transform 1 0 13156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_143
timestamp 0
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_7
timestamp 0
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 0
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_45
timestamp 0
transform 1 0 5244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_66
timestamp 0
transform 1 0 7176 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_72
timestamp 0
transform 1 0 7728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_80
timestamp 0
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_89
timestamp 0
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_120
timestamp 0
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_127
timestamp 0
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_35
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 0
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_65
timestamp 0
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_73
timestamp 0
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_79
timestamp 0
transform 1 0 8372 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_87
timestamp 0
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_124
timestamp 0
transform 1 0 12512 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_135
timestamp 0
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_23
timestamp 0
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_33
timestamp 0
transform 1 0 4140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_49
timestamp 0
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_57
timestamp 0
transform 1 0 6348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_80
timestamp 0
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_116
timestamp 0
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_127
timestamp 0
transform 1 0 12788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_35
timestamp 0
transform 1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_44
timestamp 0
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_95
timestamp 0
transform 1 0 9844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_104
timestamp 0
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_130
timestamp 0
transform 1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_142
timestamp 0
transform 1 0 14168 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_19
timestamp 0
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_23
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_36
timestamp 0
transform 1 0 4416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_45
timestamp 0
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_64
timestamp 0
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_76
timestamp 0
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_98
timestamp 0
transform 1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_134
timestamp 0
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_12
timestamp 0
transform 1 0 2208 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_20
timestamp 0
transform 1 0 2944 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_38
timestamp 0
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_50
timestamp 0
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_65
timestamp 0
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_73
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_88
timestamp 0
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_99
timestamp 0
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_120
timestamp 0
transform 1 0 12144 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_132
timestamp 0
transform 1 0 13248 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_144
timestamp 0
transform 1 0 14352 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_22
timestamp 0
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_73
timestamp 0
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 0
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_89
timestamp 0
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_96
timestamp 0
transform 1 0 9936 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_108
timestamp 0
transform 1 0 11040 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_120
timestamp 0
transform 1 0 12144 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 0
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_23
timestamp 0
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_28
timestamp 0
transform 1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_35
timestamp 0
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_48
timestamp 0
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_74
timestamp 0
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_82
timestamp 0
transform 1 0 8648 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_103
timestamp 0
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_120
timestamp 0
transform 1 0 12144 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_132
timestamp 0
transform 1 0 13248 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 0
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_44
timestamp 0
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_52
timestamp 0
transform 1 0 5888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_58
timestamp 0
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_63
timestamp 0
transform 1 0 6900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_69
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_79
timestamp 0
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_102
timestamp 0
transform 1 0 10488 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_117
timestamp 0
transform 1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_36
timestamp 0
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_48
timestamp 0
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_62
timestamp 0
transform 1 0 6808 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_68
timestamp 0
transform 1 0 7360 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_76
timestamp 0
transform 1 0 8096 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_103
timestamp 0
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_119
timestamp 0
transform 1 0 12052 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_131
timestamp 0
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_143
timestamp 0
transform 1 0 14260 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_40
timestamp 0
transform 1 0 4784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_48
timestamp 0
transform 1 0 5520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_63
timestamp 0
transform 1 0 6900 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_73
timestamp 0
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 0
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_96
timestamp 0
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_106
timestamp 0
transform 1 0 10856 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_113
timestamp 0
transform 1 0 11500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_125
timestamp 0
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 0
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_36
timestamp 0
transform 1 0 4416 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_40
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_52
timestamp 0
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_78
timestamp 0
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_90
timestamp 0
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_102
timestamp 0
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_145
timestamp 0
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_47
timestamp 0
transform 1 0 5428 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_59
timestamp 0
transform 1 0 6532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 0
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_95
timestamp 0
transform 1 0 9844 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_103
timestamp 0
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_113
timestamp 0
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_125
timestamp 0
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 0
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_9
timestamp 0
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_21
timestamp 0
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_25
timestamp 0
transform 1 0 3404 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_45
timestamp 0
transform 1 0 5244 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_64
timestamp 0
transform 1 0 6992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_79
timestamp 0
transform 1 0 8372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_100
timestamp 0
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_145
timestamp 0
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_57
timestamp 0
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_69
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_41
timestamp 0
transform 1 0 4876 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_46
timestamp 0
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 0
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_65
timestamp 0
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_79
timestamp 0
transform 1 0 8372 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_86
timestamp 0
transform 1 0 9016 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_98
timestamp 0
transform 1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_107
timestamp 0
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_135
timestamp 0
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_33
timestamp 0
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_106
timestamp 0
transform 1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_118
timestamp 0
transform 1 0 11960 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_130
timestamp 0
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 0
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_9
timestamp 0
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_21
timestamp 0
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_33
timestamp 0
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_45
timestamp 0
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 0
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_72
timestamp 0
transform 1 0 7728 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_84
timestamp 0
transform 1 0 8832 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_96
timestamp 0
transform 1 0 9936 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_108
timestamp 0
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_12
timestamp 0
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_16
timestamp 0
transform 1 0 2576 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_20
timestamp 0
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 0
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_57
timestamp 0
transform 1 0 6348 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_72
timestamp 0
transform 1 0 7728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_90
timestamp 0
transform 1 0 9384 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_102
timestamp 0
transform 1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_110
timestamp 0
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_113
timestamp 0
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 0
transform -1 0 14628 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 0
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 0
transform -1 0 13156 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input6
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 0
transform -1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 0
transform -1 0 13984 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input13
timestamp 0
transform 1 0 11684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input14
timestamp 0
transform -1 0 13984 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 0
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 0
transform -1 0 9384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 0
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 0
transform 1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 0
transform -1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap31
timestamp 0
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 0
transform -1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 0
transform 1 0 14076 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 0
transform 1 0 14076 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 0
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 0
transform -1 0 7728 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 0
transform -1 0 8832 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 0
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 0
transform -1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output30
timestamp 0
transform 1 0 13800 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 14904 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 14904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 14904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 14904 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 14904 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 14904 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 14904 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
<< labels >>
rlabel metal1 s 8004 15232 8004 15232 4 VGND
rlabel metal1 s 8004 15776 8004 15776 4 VPWR
rlabel metal1 s 11914 6256 11914 6256 4 _000_
rlabel metal2 s 7406 13396 7406 13396 4 _001_
rlabel metal1 s 7958 13770 7958 13770 4 _002_
rlabel metal1 s 5658 10064 5658 10064 4 _003_
rlabel metal2 s 7498 9860 7498 9860 4 _004_
rlabel metal1 s 6900 9418 6900 9418 4 _005_
rlabel metal1 s 7820 9350 7820 9350 4 _006_
rlabel metal1 s 7314 11050 7314 11050 4 _007_
rlabel metal1 s 8326 10166 8326 10166 4 _008_
rlabel metal1 s 8832 6766 8832 6766 4 _009_
rlabel metal1 s 8464 11050 8464 11050 4 _010_
rlabel metal1 s 7958 9690 7958 9690 4 _011_
rlabel metal1 s 8096 9418 8096 9418 4 _012_
rlabel metal1 s 11040 10234 11040 10234 4 _013_
rlabel metal2 s 11178 10948 11178 10948 4 _014_
rlabel metal1 s 10856 11322 10856 11322 4 _015_
rlabel metal1 s 9338 12886 9338 12886 4 _016_
rlabel metal1 s 9012 12954 9012 12954 4 _017_
rlabel metal1 s 9844 13226 9844 13226 4 _018_
rlabel metal1 s 9522 11322 9522 11322 4 _019_
rlabel metal1 s 9706 11866 9706 11866 4 _020_
rlabel metal2 s 9246 9860 9246 9860 4 _021_
rlabel metal2 s 9890 10948 9890 10948 4 _022_
rlabel metal1 s 10626 11832 10626 11832 4 _023_
rlabel metal1 s 11132 11730 11132 11730 4 _024_
rlabel metal1 s 10074 7922 10074 7922 4 _025_
rlabel metal1 s 10350 9607 10350 9607 4 _026_
rlabel metal1 s 10258 8432 10258 8432 4 _027_
rlabel metal1 s 9844 9622 9844 9622 4 _028_
rlabel metal1 s 9246 8568 9246 8568 4 _029_
rlabel metal1 s 9292 8058 9292 8058 4 _030_
rlabel metal1 s 8050 7446 8050 7446 4 _031_
rlabel metal1 s 13110 6732 13110 6732 4 _032_
rlabel metal1 s 8602 7480 8602 7480 4 _033_
rlabel metal1 s 11224 8942 11224 8942 4 _034_
rlabel metal2 s 11546 9248 11546 9248 4 _035_
rlabel metal1 s 11546 7242 11546 7242 4 _036_
rlabel metal1 s 11684 8602 11684 8602 4 _037_
rlabel metal1 s 9614 8500 9614 8500 4 _038_
rlabel metal1 s 9798 6766 9798 6766 4 _039_
rlabel metal1 s 9522 6732 9522 6732 4 _040_
rlabel metal1 s 9292 6834 9292 6834 4 _041_
rlabel metal1 s 12834 6834 12834 6834 4 _042_
rlabel metal1 s 11822 6732 11822 6732 4 _043_
rlabel metal1 s 11408 4794 11408 4794 4 _044_
rlabel metal1 s 10902 5882 10902 5882 4 _045_
rlabel metal1 s 11730 6800 11730 6800 4 _046_
rlabel metal2 s 10994 6596 10994 6596 4 _047_
rlabel metal2 s 10534 4828 10534 4828 4 _048_
rlabel metal1 s 10672 6426 10672 6426 4 _049_
rlabel metal1 s 11500 6766 11500 6766 4 _050_
rlabel metal1 s 10166 6834 10166 6834 4 _051_
rlabel metal1 s 8326 4012 8326 4012 4 _052_
rlabel metal1 s 12581 4998 12581 4998 4 _053_
rlabel metal1 s 7958 5236 7958 5236 4 _054_
rlabel metal1 s 8142 4692 8142 4692 4 _055_
rlabel metal1 s 8694 3026 8694 3026 4 _056_
rlabel metal2 s 9246 4250 9246 4250 4 _057_
rlabel metal1 s 9706 5100 9706 5100 4 _058_
rlabel metal1 s 9798 5202 9798 5202 4 _059_
rlabel metal3 s 9154 4556 9154 4556 4 _060_
rlabel metal1 s 9522 3162 9522 3162 4 _061_
rlabel metal1 s 9936 3706 9936 3706 4 _062_
rlabel metal1 s 10212 3706 10212 3706 4 _063_
rlabel metal1 s 10258 4148 10258 4148 4 _064_
rlabel metal1 s 9568 4046 9568 4046 4 _065_
rlabel metal1 s 8648 4250 8648 4250 4 _066_
rlabel metal1 s 7084 2958 7084 2958 4 _067_
rlabel metal1 s 5290 3094 5290 3094 4 _068_
rlabel metal1 s 5474 3094 5474 3094 4 _069_
rlabel metal1 s 5842 2992 5842 2992 4 _070_
rlabel metal1 s 7774 2618 7774 2618 4 _071_
rlabel metal1 s 7958 2992 7958 2992 4 _072_
rlabel metal1 s 5842 2856 5842 2856 4 _073_
rlabel metal1 s 5244 5134 5244 5134 4 _074_
rlabel metal1 s 4692 4114 4692 4114 4 _075_
rlabel metal1 s 5750 3060 5750 3060 4 _076_
rlabel metal1 s 5290 2890 5290 2890 4 _077_
rlabel metal1 s 6072 3162 6072 3162 4 _078_
rlabel metal2 s 7590 10234 7590 10234 4 _079_
rlabel metal1 s 8694 8942 8694 8942 4 _080_
rlabel metal1 s 6532 4794 6532 4794 4 _081_
rlabel metal1 s 4002 7888 4002 7888 4 _082_
rlabel metal1 s 6762 7854 6762 7854 4 _083_
rlabel metal1 s 3634 6698 3634 6698 4 _084_
rlabel metal2 s 11730 10302 11730 10302 4 _085_
rlabel metal2 s 6578 8296 6578 8296 4 _086_
rlabel metal1 s 6486 7888 6486 7888 4 _087_
rlabel metal1 s 4600 8874 4600 8874 4 _088_
rlabel metal1 s 5428 8602 5428 8602 4 _089_
rlabel metal1 s 6348 8466 6348 8466 4 _090_
rlabel metal1 s 4508 6970 4508 6970 4 _091_
rlabel metal1 s 6486 9520 6486 9520 4 _092_
rlabel metal1 s 10166 9486 10166 9486 4 _093_
rlabel metal1 s 11132 6766 11132 6766 4 _094_
rlabel metal1 s 4324 8602 4324 8602 4 _095_
rlabel metal1 s 6256 8398 6256 8398 4 _096_
rlabel metal1 s 12512 5202 12512 5202 4 _097_
rlabel metal1 s 12466 5304 12466 5304 4 _098_
rlabel metal2 s 12650 6596 12650 6596 4 _099_
rlabel metal1 s 10971 7786 10971 7786 4 _100_
rlabel metal1 s 6026 5338 6026 5338 4 _101_
rlabel metal1 s 5612 4114 5612 4114 4 _102_
rlabel metal1 s 7544 4794 7544 4794 4 _103_
rlabel metal2 s 6394 3978 6394 3978 4 _104_
rlabel metal1 s 10074 3162 10074 3162 4 _105_
rlabel metal1 s 10028 4590 10028 4590 4 _106_
rlabel metal1 s 8142 6256 8142 6256 4 _107_
rlabel metal2 s 9890 13090 9890 13090 4 _108_
rlabel metal1 s 7590 10710 7590 10710 4 _109_
rlabel metal1 s 4876 12818 4876 12818 4 _110_
rlabel metal1 s 4922 12886 4922 12886 4 _111_
rlabel metal1 s 4692 11866 4692 11866 4 _112_
rlabel metal1 s 4830 12648 4830 12648 4 _113_
rlabel metal1 s 10626 13294 10626 13294 4 _114_
rlabel metal1 s 10304 12954 10304 12954 4 _115_
rlabel metal1 s 8602 13396 8602 13396 4 _116_
rlabel metal1 s 8004 7922 8004 7922 4 _117_
rlabel metal1 s 6670 5644 6670 5644 4 _118_
rlabel metal1 s 9982 2482 9982 2482 4 _119_
rlabel metal1 s 13156 6426 13156 6426 4 _120_
rlabel metal2 s 13202 4046 13202 4046 4 _121_
rlabel metal1 s 11224 3162 11224 3162 4 _122_
rlabel metal1 s 8418 2482 8418 2482 4 _123_
rlabel metal2 s 7866 4692 7866 4692 4 _124_
rlabel metal1 s 6210 5746 6210 5746 4 _125_
rlabel metal1 s 5382 13362 5382 13362 4 _126_
rlabel metal1 s 6049 12954 6049 12954 4 _127_
rlabel metal1 s 8372 12682 8372 12682 4 _128_
rlabel metal1 s 6578 6222 6578 6222 4 _129_
rlabel metal2 s 7038 6086 7038 6086 4 _130_
rlabel metal1 s 7130 6324 7130 6324 4 _131_
rlabel metal1 s 6808 6290 6808 6290 4 _132_
rlabel metal1 s 7360 6426 7360 6426 4 _133_
rlabel metal1 s 6670 8874 6670 8874 4 _134_
rlabel metal2 s 5934 12002 5934 12002 4 _135_
rlabel metal1 s 5980 13362 5980 13362 4 _136_
rlabel metal1 s 7452 8602 7452 8602 4 _137_
rlabel metal1 s 5842 11866 5842 11866 4 _138_
rlabel metal1 s 6486 11730 6486 11730 4 _139_
rlabel metal1 s 6532 11322 6532 11322 4 _140_
rlabel metal1 s 4462 10642 4462 10642 4 _141_
rlabel metal1 s 7774 3672 7774 3672 4 _142_
rlabel metal1 s 3910 9690 3910 9690 4 _143_
rlabel metal1 s 5796 9894 5796 9894 4 _144_
rlabel metal1 s 5750 11696 5750 11696 4 _145_
rlabel metal1 s 3634 5678 3634 5678 4 _146_
rlabel metal1 s 11454 10642 11454 10642 4 _147_
rlabel metal1 s 4738 10778 4738 10778 4 _148_
rlabel metal1 s 5382 11322 5382 11322 4 _149_
rlabel metal1 s 14766 11118 14766 11118 4 a[0]
rlabel metal2 s 3910 1027 3910 1027 4 a[1]
rlabel metal3 s 1050 13668 1050 13668 4 a[2]
rlabel metal3 s 820 2108 820 2108 4 a[3]
rlabel metal2 s 12926 1588 12926 1588 4 a[4]
rlabel metal3 s 1096 6868 1096 6868 4 a[5]
rlabel metal3 s 820 4148 820 4148 4 a[6]
rlabel metal1 s 14720 6290 14720 6290 4 a[7]
rlabel metal2 s 4554 17011 4554 17011 4 b[0]
rlabel metal2 s 46 1588 46 1588 4 b[1]
rlabel metal1 s 13892 15402 13892 15402 4 b[2]
rlabel metal1 s 14720 15470 14720 15470 4 b[3]
rlabel metal1 s 11730 15470 11730 15470 4 b[4]
rlabel metal1 s 13846 2448 13846 2448 4 b[5]
rlabel metal2 s 10994 1588 10994 1588 4 b[6]
rlabel metal1 s 1012 15470 1012 15470 4 b[7]
rlabel metal2 s 15502 1554 15502 1554 4 carry
rlabel metal1 s 5290 13498 5290 13498 4 net1
rlabel metal1 s 2208 2618 2208 2618 4 net10
rlabel metal1 s 10396 13294 10396 13294 4 net11
rlabel metal1 s 13570 12818 13570 12818 4 net12
rlabel metal1 s 13110 5032 13110 5032 4 net13
rlabel metal1 s 12512 2482 12512 2482 4 net14
rlabel metal2 s 11086 2822 11086 2822 4 net15
rlabel metal2 s 2162 10540 2162 10540 4 net16
rlabel metal1 s 8970 15334 8970 15334 4 net17
rlabel metal1 s 2714 2618 2714 2618 4 net18
rlabel metal1 s 2944 7854 2944 7854 4 net19
rlabel metal1 s 3956 10574 3956 10574 4 net2
rlabel metal1 s 14122 4794 14122 4794 4 net20
rlabel metal1 s 14076 2414 14076 2414 4 net21
rlabel metal1 s 7360 9010 7360 9010 4 net22
rlabel metal1 s 14076 13906 14076 13906 4 net23
rlabel metal1 s 14030 14994 14030 14994 4 net24
rlabel metal1 s 7544 9078 7544 9078 4 net25
rlabel metal1 s 7636 15402 7636 15402 4 net26
rlabel metal1 s 9246 2346 9246 2346 4 net27
rlabel metal1 s 1794 8976 1794 8976 4 net28
rlabel metal1 s 3772 15402 3772 15402 4 net29
rlabel metal1 s 10810 13396 10810 13396 4 net3
rlabel metal1 s 13938 8534 13938 8534 4 net30
rlabel metal1 s 9338 8432 9338 8432 4 net31
rlabel metal1 s 4002 2550 4002 2550 4 net4
rlabel metal2 s 12834 6052 12834 6052 4 net5
rlabel metal1 s 2415 7446 2415 7446 4 net6
rlabel metal2 s 4830 4114 4830 4114 4 net7
rlabel metal1 s 6164 5202 6164 5202 4 net8
rlabel metal1 s 4692 13498 4692 13498 4 net9
rlabel metal1 s 9200 15470 9200 15470 4 opcode[0]
rlabel metal2 s 1978 1588 1978 1588 4 opcode[1]
rlabel metal2 s 2622 17011 2622 17011 4 opcode[2]
rlabel metal1 s 14766 4590 14766 4590 4 opcode[3]
rlabel metal2 s 6486 1520 6486 1520 4 result[0]
rlabel metal1 s 14674 13838 14674 13838 4 result[1]
rlabel metal1 s 14674 15130 14674 15130 4 result[2]
rlabel metal3 s 820 11628 820 11628 4 result[3]
rlabel metal2 s 7130 17011 7130 17011 4 result[4]
rlabel metal2 s 8418 1520 8418 1520 4 result[5]
rlabel metal3 s 820 8908 820 8908 4 result[6]
rlabel metal3 s 820 16388 820 16388 4 result[7]
rlabel metal2 s 14490 8721 14490 8721 4 zero
flabel metal4 s 4868 2128 5188 15824 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 15346 14952 15666 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5346 14952 5666 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 14208 2128 14528 15824 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4208 2128 4528 15824 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 15289 10888 16089 11008 0 FreeSans 600 0 0 0 a[0]
port 3 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 a[1]
port 4 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 a[2]
port 5 nsew
flabel metal3 s 0 2048 800 2168 0 FreeSans 600 0 0 0 a[3]
port 6 nsew
flabel metal2 s 12898 0 12954 800 0 FreeSans 280 90 0 0 a[4]
port 7 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 a[5]
port 8 nsew
flabel metal3 s 0 4088 800 4208 0 FreeSans 600 0 0 0 a[6]
port 9 nsew
flabel metal3 s 15289 6128 16089 6248 0 FreeSans 600 0 0 0 a[7]
port 10 nsew
flabel metal2 s 4526 17433 4582 18233 0 FreeSans 280 90 0 0 b[0]
port 11 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 b[1]
port 12 nsew
flabel metal2 s 13542 17433 13598 18233 0 FreeSans 280 90 0 0 b[2]
port 13 nsew
flabel metal2 s 15474 17433 15530 18233 0 FreeSans 280 90 0 0 b[3]
port 14 nsew
flabel metal2 s 11610 17433 11666 18233 0 FreeSans 280 90 0 0 b[4]
port 15 nsew
flabel metal3 s 15289 1368 16089 1488 0 FreeSans 600 0 0 0 b[5]
port 16 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 b[6]
port 17 nsew
flabel metal2 s 18 17433 74 18233 0 FreeSans 280 90 0 0 b[7]
port 18 nsew
flabel metal2 s 15474 0 15530 800 0 FreeSans 280 90 0 0 carry
port 19 nsew
flabel metal2 s 9034 17433 9090 18233 0 FreeSans 280 90 0 0 opcode[0]
port 20 nsew
flabel metal2 s 1950 0 2006 800 0 FreeSans 280 90 0 0 opcode[1]
port 21 nsew
flabel metal2 s 2594 17433 2650 18233 0 FreeSans 280 90 0 0 opcode[2]
port 22 nsew
flabel metal3 s 15289 4088 16089 4208 0 FreeSans 600 0 0 0 opcode[3]
port 23 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 result[0]
port 24 nsew
flabel metal3 s 15289 13608 16089 13728 0 FreeSans 600 0 0 0 result[1]
port 25 nsew
flabel metal3 s 15289 15648 16089 15768 0 FreeSans 600 0 0 0 result[2]
port 26 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 result[3]
port 27 nsew
flabel metal2 s 7102 17433 7158 18233 0 FreeSans 280 90 0 0 result[4]
port 28 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 result[5]
port 29 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 result[6]
port 30 nsew
flabel metal3 s 0 16328 800 16448 0 FreeSans 600 0 0 0 result[7]
port 31 nsew
flabel metal3 s 15289 8848 16089 8968 0 FreeSans 600 0 0 0 zero
port 32 nsew
<< properties >>
string FIXED_BBOX 0 0 16089 18233
<< end >>
